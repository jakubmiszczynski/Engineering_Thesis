** sch_path: /home/kuba/project/SKY130_OpAmp/06_ParasiticsSim/opamp_cascode_ac_ochoa_mc.sch
**.subckt opamp_cascode_ac_ochoa_mc
V2 Vout net1 DC=0 AC={B}
.save i(v2)
C1 Vout GND 1p m=1
C2 VoutQ GND 1p m=1
V1 net2 net1 DC=0 AC={1-B}
.save i(v1)
B1 net1 GND v=V(VoutQ)
I0 IBIAS GND 45u
x1 Vp net2 VCC GND Vout VB_A VB_B IBIAS opamp_cascode
x2 Vp VoutQ VCC GND VoutQ VB_A VB_B IBIAS opamp_cascode
**** begin user architecture code


Vsupply VCC GND 1.8
VbiasA VB_A GND 0.2
VbiasB VB_B GND 1.1
Vin Vp GND 0.9
.param B=0
.include ../opamp_cascode.spice
.control
  set wr_vecnames
  set wr_singlescale
  let mc_runs=3
  let run=1
  set curplot=new
  set final=$curplot
  setplot $final
  dowhile run <= mc_runs
    alterparam B=0
    reset
    ac dec 10 1 1G
    alterparam B=1
    reset
    ac dec 10 1 1G
    let ixf = 2*run-1
    let ixs = 2*run
    let frequency = ac{$&ixf}.frequency
    let T = (ac{$&ixf}.i(V2) + ac{$&ixs}.i(V1)) / (ac{$&ixf}.i(V1) + ac{$&ixs}.i(V2))
    let mag = db(T)
    let phase = 180*cph(T)/pi
    set dt = $curplot
    setplot $final
    let mag{$&run}={$dt}.mag
    let phase{$&run}={$dt}.phase
    setplot $dt
    let run = run + 1
  end
  setplot $final
  plot all vs ac1.frequency xlog
.endc



.param mc_mm_switch=1
.param mc_pr_switch=0
.include ~/.volare/sky130A/libs.tech/ngspice/corners/ss.spice
.include ~/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include ~/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include ~/.volare/sky130A/libs.tech/ngspice/corners/ss/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
