* NGSPICE file created from opamp_cascode.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_SCE452 a_n158_n125# a_n100_n213# a_100_n125# VSUBS
X0 a_100_n125# a_n100_n213# a_n158_n125# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
.ends

.subckt sky130_fd_pr__pfet_01v8_ZLZ7XS w_n1594_n600# a_n1500_n597# a_1500_n500# a_n1558_n500#
X0 a_1500_n500# a_n1500_n597# a_n1558_n500# w_n1594_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__pfet_01v8_7DHACV w_n112_636# a_n33_n5541# a_n33_n8013# a_n76_736#
+ w_n112_1872# w_n112_4344# a_18_n500# a_18_n2972# a_18_n5444# a_n76_n1736# a_n33_3111#
+ a_n76_n4208# a_18_3208# a_n76_n7916# a_n33_n1833# a_18_6916# a_n76_5680# w_n112_n3072#
+ a_n33_n4305# a_n33_5583# a_n76_8152# w_n112_n6780# a_n33_8055# a_n33_n3069# a_n33_639#
+ w_n112_n9252# w_n112_3108# w_n112_6816# a_n33_n6777# a_n33_n597# a_n33_n9249# a_18_n1736#
+ a_18_n4208# a_18_n7916# a_n76_1972# a_n33_1875# w_n112_n600# a_n76_n6680# a_18_736#
+ a_n76_4444# a_18_5680# a_n33_4347# w_n112_n5544# a_n76_n9152# a_18_8152# w_n112_n8016#
+ a_n76_n500# w_n112_5580# w_n112_8052# a_18_n6680# a_n76_n2972# a_18_1972# a_n76_3208#
+ a_n76_n5444# a_18_4444# a_n76_6916# w_n112_n1836# a_18_n9152# a_n33_6819# w_n112_n4308#
X0 a_18_3208# a_n33_3111# a_n76_3208# w_n112_3108# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1 a_18_n6680# a_n33_n6777# a_n76_n6680# w_n112_n6780# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X2 a_18_n500# a_n33_n597# a_n76_n500# w_n112_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X3 a_18_n9152# a_n33_n9249# a_n76_n9152# w_n112_n9252# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X4 a_18_736# a_n33_639# a_n76_736# w_n112_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X5 a_18_n2972# a_n33_n3069# a_n76_n2972# w_n112_n3072# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X6 a_18_n7916# a_n33_n8013# a_n76_n7916# w_n112_n8016# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X7 a_18_5680# a_n33_5583# a_n76_5680# w_n112_5580# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X8 a_18_n5444# a_n33_n5541# a_n76_n5444# w_n112_n5544# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X9 a_18_8152# a_n33_8055# a_n76_8152# w_n112_8052# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X10 a_18_n1736# a_n33_n1833# a_n76_n1736# w_n112_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X11 a_18_6916# a_n33_6819# a_n76_6916# w_n112_6816# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X12 a_18_1972# a_n33_1875# a_n76_1972# w_n112_1872# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X13 a_18_n4208# a_n33_n4305# a_n76_n4208# w_n112_n4308# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X14 a_18_4444# a_n33_4347# a_n76_4444# w_n112_4344# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__nfet_01v8_MHE452 a_n158_n359# a_n100_957# a_100_n1295# a_n158_577#
+ a_n100_21# a_100_109# a_n100_n915# a_100_n827# a_n100_489# a_100_1045# a_n158_n1295#
+ a_n158_n827# a_100_577# a_n158_1045# a_n100_n447# a_n158_109# a_100_n359# a_n100_n1383#
+ VSUBS
X0 a_100_n827# a_n100_n915# a_n158_n827# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X1 a_100_n359# a_n100_n447# a_n158_n359# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X2 a_100_577# a_n100_489# a_n158_577# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X3 a_100_1045# a_n100_957# a_n158_1045# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X4 a_100_n1295# a_n100_n1383# a_n158_n1295# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X5 a_100_109# a_n100_21# a_n158_109# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
.ends

.subckt sky130_fd_pr__pfet_01v8_P2UXFR a_n300_n1215# w_n394_n1218# a_n358_n1118# a_n300_21#
+ a_300_118# w_n394_18# a_300_n1118# a_n358_118#
X0 a_300_118# a_n300_21# a_n358_118# w_n394_18# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X1 a_300_n1118# a_n300_n1215# a_n358_n1118# w_n394_n1218# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__nfet_01v8_VT3ZQW a_n158_n125# a_n100_n213# a_100_n125# VSUBS
X0 a_100_n125# a_n100_n213# a_n158_n125# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
.ends

.subckt sky130_fd_pr__pfet_01v8_RRUZAE a_n358_n2972# a_n300_n1833# a_n300_n3069# w_n394_n1836#
+ w_n394_1872# a_n358_n1736# a_300_736# a_300_1972# a_300_n2972# w_n394_636# w_n394_n3072#
+ a_n300_n597# a_300_n500# a_n300_639# a_n358_1972# a_n300_1875# w_n394_n600# a_300_n1736#
+ a_n358_n500# a_n358_736#
X0 a_300_n500# a_n300_n597# a_n358_n500# w_n394_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X1 a_300_736# a_n300_639# a_n358_736# w_n394_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X2 a_300_n2972# a_n300_n3069# a_n358_n2972# w_n394_n3072# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X3 a_300_1972# a_n300_1875# a_n358_1972# w_n394_1872# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X4 a_300_n1736# a_n300_n1833# a_n358_n1736# w_n394_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__pfet_01v8_F76D73 a_n1558_11242# a_n1558_n14714# a_n1500_n43239#
+ w_n1594_n3690# a_n1500_n11103# a_n1558_50794# a_1500_n23366# a_n1500_n50655# w_n1594_n56838#
+ w_n1594_n24702# a_1500_n30782# a_n1500_3729# a_n1558_n60446# w_n1594_12378# a_1500_n8534#
+ a_n1558_14950# a_1500_n19658# a_n1500_n14811# a_n1500_n46947# w_n1594_9906# w_n1594_n6162#
+ a_1500_22366# a_n1500_22269# a_n1558_53266# a_n1558_n56738# a_n1558_n24602# a_n1558_21130#
+ a_n1500_n53127# w_n1594_n13578# a_n1558_60682# a_1500_n33254# a_n1500_n60543# w_n1594_n20994#
+ a_1500_n40670# a_1500_18658# a_n1558_49558# a_n1558_17422# w_n1594_22266# a_n1500_n49419#
+ w_n1594_n9870# a_n1500_25977# a_n1558_56974# a_n1500_n56835# a_1500_n29546# a_n1558_n3590#
+ a_1500_n36962# a_n1500_9909# a_n1558_n13478# a_1500_32254# a_n1500_32157# a_n1558_n20894#
+ w_n1594_18558# w_n1594_n23466# a_1500_n43142# w_n1594_n30882# w_n1594_25974# a_n1500_n2451#
+ a_1500_28546# a_1500_n7298# a_n1500_28449# a_n1558_59446# a_n1558_27310# a_n1500_n13575#
+ a_n1500_n59307# w_n1594_32154# w_n1594_n19758# a_1500_35962# a_n1558_n6062# a_n1500_35865#
+ a_1500_n39434# a_n1500_n20991# a_1500_n46850# a_n1558_n23366# a_1500_42142# a_n1500_42045#
+ a_n1558_n30782# w_n1594_n33354# w_n1594_28446# a_1500_n53030# w_n1594_35862# w_n1594_n40770#
+ a_n1558_n9770# w_n1594_18# a_n1558_16186# a_n1500_21# a_n1558_n19658# a_n1500_n16047#
+ a_1500_38434# a_n1500_38337# a_n1500_n55599# a_n1500_n23463# w_n1594_n29646# a_1500_45850#
+ w_n1594_42042# a_n1500_45753# a_n1558_40906# a_1500_n49322# a_n1558_n33254# a_1500_52030#
+ a_n1500_n8631# a_n1558_n40670# a_n1558_19894# w_n1594_38334# w_n1594_n43242# a_n1500_n19755#
+ w_n1594_45750# a_n1558_26074# a_n1558_n29546# a_1500_48322# a_n1500_48225# a_1500_n38198#
+ a_n1558_33490# a_n1558_n36962# a_n1500_n33351# w_n1594_n39534# a_n1500_55641# a_1500_n59210#
+ w_n1594_n46950# a_n1558_n43142# a_n1558_29782# w_n1594_n53130# a_n1500_n29643# w_n1594_48222#
+ a_1500_37198# a_n1558_n39434# a_1500_58210# a_n1500_58113# a_n1500_12381# a_1500_n1118#
+ a_1500_n48086# a_n1558_n46850# w_n1594_n49422# a_n1500_n7395# a_n1558_n53030# w_n1594_37098#
+ a_n1558_39670# a_n1500_n39531# w_n1594_58110# a_1500_n4826# a_1500_47086# a_n1558_10006#
+ a_n1558_n49322# w_n1594_n2454# w_n1594_n38298# a_1500_2590# w_n1594_2490# w_n1594_n59310#
+ a_n1500_6201# a_n1500_18561# a_n1558_13714# a_n1558_2590# a_1500_n25838# a_n1558_n38198#
+ a_1500_5062# a_1500_118# a_n1558_n59210# w_n1594_n48186# w_n1594_n16050# a_1500_n32018#
+ a_n1500_2493# a_1500_24838# a_n1558_5062# a_n1500_n38295# w_n1594_n8634# a_1500_8770#
+ a_n1558_55738# a_n1558_23602# a_n1558_n2354# w_n1594_8670# a_1500_n35726# a_n1558_n48086#
+ a_1500_31018# w_n1594_n58074# w_n1594_24738# a_n1558_8770# a_n1500_n1215# a_n1558_12478#
+ a_n1500_n12339# a_n1500_n48183# a_1500_34726# a_n1500_34629# w_n1594_n25938# a_1500_n45614#
+ a_n1500_8673# w_n1594_n32118# a_n1500_n4923# w_n1594_34626# a_n1558_n8534# w_n1594_n7398#
+ a_n1558_22366# a_n1558_n25838# a_n1500_n22227# a_n1500_n58071# a_1500_44614# a_n1500_44517#
+ a_n1500_n61779# w_n1594_n35826# a_n1500_51933# a_1500_n55502# a_n1558_n32018# a_n1558_18658#
+ w_n1594_n42006# a_n1500_n18519# a_n1500_n25935# w_n1594_44514# w_n1594_51930# a_n1558_32254#
+ a_n1558_n35726# a_n1500_n32115# a_1500_54502# a_n1500_54405# a_1500_n44378# a_1500_n12242#
+ w_n1594_n45714# a_1500_n51794# a_n1500_n3687# a_n1558_28546# a_n1558_n7298# a_n1500_n28407#
+ a_n1558_35962# a_n1500_n35823# w_n1594_54402# a_1500_n15950# a_1500_43378# a_1500_11242#
+ a_n1500_11145# a_n1558_42142# a_n1558_n45614# a_1500_50794# a_n1500_n42003# a_n1500_50697#
+ a_1500_n54266# a_1500_n22130# a_n1500_n6159# w_n1594_n55602# a_1500_n61682# a_n1558_38434#
+ a_n1500_n24699# w_n1594_43278# w_n1594_11142# a_1500_14950# a_n1500_46989# a_n1558_45850#
+ a_n1500_14853# a_1500_n18422# a_n1500_n45711# w_n1594_50694# a_1500_n57974# a_n1500_n9867#
+ w_n1594_n1218# a_1500_53266# a_1500_1354# a_n1500_53169# a_1500_21130# a_n1500_21033#
+ a_n1558_n55502# a_n1558_52030# w_n1594_1254# w_n1594_n12342# w_n1594_n44478# a_1500_60682#
+ a_n1500_60585# w_n1594_14850# w_n1594_n51894# w_n1594_46986# a_1500_49558# a_1500_17422#
+ a_n1558_48322# a_n1500_17325# a_n1500_n34587# a_1500_56974# a_n1558_1354# w_n1594_53166#
+ w_n1594_21030# w_n1594_n4926# a_n1500_56877# a_n1500_24741# a_1500_n3590# a_1500_n28310#
+ w_n1594_60582# w_n1594_4962# a_n1558_n44378# a_n1558_n12242# a_n1558_n51794# w_n1594_17322#
+ w_n1594_n22230# w_n1594_n54366# w_n1594_49458# a_n1500_1257# w_n1594_n61782# w_n1594_56874#
+ a_n1558_37198# a_n1500_n37059# a_1500_59446# a_1500_27310# a_1500_7534# a_n1500_59349#
+ a_n1500_27213# a_1500_n6062# a_1500_n17186# a_n1558_58210# a_n1558_n15950# a_n1500_n44475#
+ a_n1558_n1118# w_n1594_7434# w_n1594_n18522# a_n1500_n51891# a_n1558_n54266# a_1500_n41906#
+ a_n1500_4965# a_n1558_n22130# a_n1558_n61682# w_n1594_59346# w_n1594_27210# a_n1558_7534#
+ a_1500_n9770# w_n1594_30918# a_n1558_n4826# a_1500_16186# a_n1500_16089# a_n1558_47086#
+ a_n1558_n18422# a_n1500_37101# a_n1558_n57974# a_1500_n27074# a_n1500_n54363# a_1500_40906#
+ w_n1594_n28410# a_n1500_40809# a_1500_n34490# a_n1500_7437# w_n1594_16086# a_1500_19894#
+ a_n1500_19797# w_n1594_40806# a_1500_26074# a_1500_6298# a_n1558_n28310# w_n1594_6198#
+ w_n1594_n17286# a_1500_33490# a_n1500_33393# w_n1594_19794# a_n1558_6298# a_1500_29782#
+ a_n1500_29685# a_n1558_24838# w_n1594_33390# a_n1558_n17186# a_n1558_118# a_n1558_31018#
+ w_n1594_n27174# a_n1500_43281# a_n1558_n41906# a_1500_n11006# w_n1594_29682# w_n1594_n34590#
+ a_1500_n50558# a_n1500_n17283# a_1500_39670# a_n1500_39573# a_n1558_34726# a_1500_n14714#
+ a_n1558_n27074# a_1500_10006# a_n1558_n34490# w_n1594_n37062# w_n1594_39570# a_1500_n60446#
+ a_n1500_n27171# a_1500_13714# a_n1500_13617# a_n1500_49461# a_n1558_44614# a_n1500_n30879#
+ a_1500_n56738# a_1500_n24602# w_n1594_n11106# w_n1594_n50658# w_n1594_13614# a_1500_55738#
+ a_1500_23602# a_1500_3826# a_n1500_23505# a_1500_n2354# a_1500_n13478# a_n1558_54502#
+ a_n1500_n40767# w_n1594_3726# w_n1594_n14814# a_n1500_30921# a_1500_n20894# a_n1558_n11006#
+ a_n1558_n50558# w_n1594_n60546# a_n1558_3826# w_n1594_55638# w_n1594_23502# a_1500_12478#
+ a_n1558_43378#
X0 a_1500_53266# a_n1500_53169# a_n1558_53266# w_n1594_53166# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1 a_1500_n18422# a_n1500_n18519# a_n1558_n18422# w_n1594_n18522# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X2 a_1500_n45614# a_n1500_n45711# a_n1558_n45614# w_n1594_n45714# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X3 a_1500_n43142# a_n1500_n43239# a_n1558_n43142# w_n1594_n43242# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X4 a_1500_n22130# a_n1500_n22227# a_n1558_n22130# w_n1594_n22230# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X5 a_1500_n3590# a_n1500_n3687# a_n1558_n3590# w_n1594_n3690# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X6 a_1500_35962# a_n1500_35865# a_n1558_35962# w_n1594_35862# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X7 a_1500_33490# a_n1500_33393# a_n1558_33490# w_n1594_33390# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X8 a_1500_60682# a_n1500_60585# a_n1558_60682# w_n1594_60582# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X9 a_1500_12478# a_n1500_12381# a_n1558_12478# w_n1594_12378# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X10 a_1500_38434# a_n1500_38337# a_n1558_38434# w_n1594_38334# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X11 a_1500_6298# a_n1500_6201# a_n1558_6298# w_n1594_6198# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X12 a_1500_n55502# a_n1500_n55599# a_n1558_n55502# w_n1594_n55602# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X13 a_1500_n32018# a_n1500_n32115# a_n1558_n32018# w_n1594_n32118# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X14 a_1500_45850# a_n1500_45753# a_n1558_45850# w_n1594_45750# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X15 a_1500_24838# a_n1500_24741# a_n1558_24838# w_n1594_24738# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X16 a_1500_n38198# a_n1500_n38295# a_n1558_n38198# w_n1594_n38298# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X17 a_1500_22366# a_n1500_22269# a_n1558_22366# w_n1594_22266# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X18 a_1500_48322# a_n1500_48225# a_n1558_48322# w_n1594_48222# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X19 a_1500_n14714# a_n1500_n14811# a_n1558_n14714# w_n1594_n14814# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X20 a_1500_n41906# a_n1500_n42003# a_n1558_n41906# w_n1594_n42006# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X21 a_1500_n12242# a_n1500_n12339# a_n1558_n12242# w_n1594_n12342# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X22 a_1500_34726# a_n1500_34629# a_n1558_34726# w_n1594_34626# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X23 a_1500_32254# a_n1500_32157# a_n1558_32254# w_n1594_32154# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X24 a_1500_n48086# a_n1500_n48183# a_n1558_n48086# w_n1594_n48186# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X25 a_1500_58210# a_n1500_58113# a_n1558_58210# w_n1594_58110# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X26 a_1500_n24602# a_n1500_n24699# a_n1558_n24602# w_n1594_n24702# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X27 a_1500_14950# a_n1500_14853# a_n1558_14950# w_n1594_14850# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X28 a_1500_n8534# a_n1500_n8631# a_n1558_n8534# w_n1594_n8634# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X29 a_1500_n57974# a_n1500_n58071# a_n1558_n57974# w_n1594_n58074# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X30 a_1500_n6062# a_n1500_n6159# a_n1558_n6062# w_n1594_n6162# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X31 a_1500_n34490# a_n1500_n34587# a_n1558_n34490# w_n1594_n34590# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X32 a_1500_17422# a_n1500_17325# a_n1558_17422# w_n1594_17322# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X33 a_1500_44614# a_n1500_44517# a_n1558_44614# w_n1594_44514# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X34 a_1500_42142# a_n1500_42045# a_n1558_42142# w_n1594_42042# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X35 a_1500_8770# a_n1500_8673# a_n1558_8770# w_n1594_8670# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X36 a_1500_n11006# a_n1500_n11103# a_n1558_n11006# w_n1594_n11106# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X37 a_1500_n19658# a_n1500_n19755# a_n1558_n19658# w_n1594_n19758# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X38 a_1500_n46850# a_n1500_n46947# a_n1558_n46850# w_n1594_n46950# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X39 a_1500_n17186# a_n1500_n17283# a_n1558_n17186# w_n1594_n17286# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X40 a_1500_27310# a_n1500_27213# a_n1558_27310# w_n1594_27210# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X41 a_1500_n44378# a_n1500_n44475# a_n1558_n44378# w_n1594_n44478# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X42 a_1500_54502# a_n1500_54405# a_n1558_54502# w_n1594_54402# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X43 a_1500_52030# a_n1500_51933# a_n1558_52030# w_n1594_51930# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X44 a_1500_31018# a_n1500_30921# a_n1558_31018# w_n1594_30918# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X45 a_1500_n4826# a_n1500_n4923# a_n1558_n4826# w_n1594_n4926# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X46 a_1500_37198# a_n1500_37101# a_n1558_37198# w_n1594_37098# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X47 a_1500_n2354# a_n1500_n2451# a_n1558_n2354# w_n1594_n2454# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X48 a_1500_n51794# a_n1500_n51891# a_n1558_n51794# w_n1594_n51894# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X49 a_1500_n29546# a_n1500_n29643# a_n1558_n29546# w_n1594_n29646# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X50 a_1500_13714# a_n1500_13617# a_n1558_13714# w_n1594_13614# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X51 a_1500_n56738# a_n1500_n56835# a_n1558_n56738# w_n1594_n56838# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X52 a_1500_11242# a_n1500_11145# a_n1558_11242# w_n1594_11142# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X53 a_1500_40906# a_n1500_40809# a_n1558_40906# w_n1594_40806# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X54 a_1500_n27074# a_n1500_n27171# a_n1558_n27074# w_n1594_n27174# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X55 a_1500_n54266# a_n1500_n54363# a_n1558_n54266# w_n1594_n54366# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X56 a_1500_19894# a_n1500_19797# a_n1558_19894# w_n1594_19794# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X57 a_1500_2590# a_n1500_2493# a_n1558_2590# w_n1594_2490# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X58 a_1500_n59210# a_n1500_n59307# a_n1558_n59210# w_n1594_n59310# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X59 a_1500_7534# a_n1500_7437# a_n1558_7534# w_n1594_7434# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X60 a_1500_49558# a_n1500_49461# a_n1558_49558# w_n1594_49458# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X61 a_1500_n36962# a_n1500_n37059# a_n1558_n36962# w_n1594_n37062# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X62 a_1500_5062# a_n1500_4965# a_n1558_5062# w_n1594_4962# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X63 a_1500_47086# a_n1500_46989# a_n1558_47086# w_n1594_46986# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X64 a_1500_n15950# a_n1500_n16047# a_n1558_n15950# w_n1594_n16050# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X65 a_1500_n61682# a_n1500_n61779# a_n1558_n61682# w_n1594_n61782# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X66 a_1500_n13478# a_n1500_n13575# a_n1558_n13478# w_n1594_n13578# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X67 a_1500_23602# a_n1500_23505# a_n1558_23602# w_n1594_23502# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X68 a_1500_n40670# a_n1500_n40767# a_n1558_n40670# w_n1594_n40770# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X69 a_1500_n39434# a_n1500_n39531# a_n1558_n39434# w_n1594_n39534# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X70 a_1500_21130# a_n1500_21033# a_n1558_21130# w_n1594_21030# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X71 a_1500_29782# a_n1500_29685# a_n1558_29782# w_n1594_29682# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X72 a_1500_56974# a_n1500_56877# a_n1558_56974# w_n1594_56874# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X73 a_1500_59446# a_n1500_59349# a_n1558_59446# w_n1594_59346# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X74 a_1500_n20894# a_n1500_n20991# a_n1558_n20894# w_n1594_n20994# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X75 a_1500_n25838# a_n1500_n25935# a_n1558_n25838# w_n1594_n25938# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X76 a_1500_n23366# a_n1500_n23463# a_n1558_n23366# w_n1594_n23466# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X77 a_1500_n50558# a_n1500_n50655# a_n1558_n50558# w_n1594_n50658# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X78 a_1500_n49322# a_n1500_n49419# a_n1558_n49322# w_n1594_n49422# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X79 a_1500_n1118# a_n1500_n1215# a_n1558_n1118# w_n1594_n1218# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X80 a_1500_n9770# a_n1500_n9867# a_n1558_n9770# w_n1594_n9870# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X81 a_1500_n28310# a_n1500_n28407# a_n1558_n28310# w_n1594_n28410# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X82 a_1500_n7298# a_n1500_n7395# a_n1558_n7298# w_n1594_n7398# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X83 a_1500_10006# a_n1500_9909# a_n1558_10006# w_n1594_9906# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X84 a_1500_39670# a_n1500_39573# a_n1558_39670# w_n1594_39570# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X85 a_1500_18658# a_n1500_18561# a_n1558_18658# w_n1594_18558# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X86 a_1500_n53030# a_n1500_n53127# a_n1558_n53030# w_n1594_n53130# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X87 a_1500_3826# a_n1500_3729# a_n1558_3826# w_n1594_3726# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X88 a_1500_16186# a_n1500_16089# a_n1558_16186# w_n1594_16086# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X89 a_1500_1354# a_n1500_1257# a_n1558_1354# w_n1594_1254# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X90 a_1500_43378# a_n1500_43281# a_n1558_43378# w_n1594_43278# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X91 a_1500_n30782# a_n1500_n30879# a_n1558_n30782# w_n1594_n30882# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X92 a_1500_118# a_n1500_21# a_n1558_118# w_n1594_18# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X93 a_1500_n35726# a_n1500_n35823# a_n1558_n35726# w_n1594_n35826# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X94 a_1500_n33254# a_n1500_n33351# a_n1558_n33254# w_n1594_n33354# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X95 a_1500_n60446# a_n1500_n60543# a_n1558_n60446# w_n1594_n60546# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X96 a_1500_50794# a_n1500_50697# a_n1558_50794# w_n1594_50694# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X97 a_1500_28546# a_n1500_28449# a_n1558_28546# w_n1594_28446# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X98 a_1500_55738# a_n1500_55641# a_n1558_55738# w_n1594_55638# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X99 a_1500_26074# a_n1500_25977# a_n1558_26074# w_n1594_25974# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__nfet_01v8_WK8VRD a_n500_9156# a_n558_n10244# a_500_n2936# a_500_n5372#
+ a_n500_n1806# a_500_718# a_n500_3066# a_n500_n4242# a_n500_630# a_n500_n6678# a_n558_1936#
+ a_n558_4372# a_n558_n9026# a_n558_n6590# a_500_n500# a_500_6808# a_n500_6720# a_500_9244#
+ a_500_3154# a_500_n7808# a_n500_n9114# a_500_n4154# a_500_n1718# a_n558_n500# a_n500_n3024#
+ a_n558_6808# a_n558_9244# a_n558_n2936# a_n558_3154# a_n500_n10332# a_n558_n5372#
+ a_n558_718# a_n500_n588# a_n500_5502# a_500_8026# a_500_5590# a_n500_7938# a_500_n9026#
+ a_n500_1848# a_500_n6590# a_n500_4284# a_n500_n5460# a_n558_n7808# a_n500_n7896#
+ a_n558_8026# a_n558_n1718# a_n558_5590# a_n558_n4154# a_500_n10244# a_500_1936#
+ a_500_4372# VSUBS
X0 a_500_n10244# a_n500_n10332# a_n558_n10244# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1 a_500_4372# a_n500_4284# a_n558_4372# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X2 a_500_n6590# a_n500_n6678# a_n558_n6590# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X3 a_500_5590# a_n500_5502# a_n558_5590# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X4 a_500_n1718# a_n500_n1806# a_n558_n1718# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X5 a_500_n2936# a_n500_n3024# a_n558_n2936# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X6 a_500_n4154# a_n500_n4242# a_n558_n4154# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X7 a_500_718# a_n500_630# a_n558_718# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X8 a_500_n5372# a_n500_n5460# a_n558_n5372# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X9 a_500_6808# a_n500_6720# a_n558_6808# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X10 a_500_8026# a_n500_7938# a_n558_8026# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X11 a_500_n500# a_n500_n588# a_n558_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X12 a_500_9244# a_n500_9156# a_n558_9244# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X13 a_500_1936# a_n500_1848# a_n558_1936# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X14 a_500_n7808# a_n500_n7896# a_n558_n7808# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X15 a_500_3154# a_n500_3066# a_n558_3154# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X16 a_500_n9026# a_n500_n9114# a_n558_n9026# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__pfet_01v8_C2U9V5 a_n300_n597# a_300_n500# w_n394_n600# a_n358_n500#
X0 a_300_n500# a_n300_n597# a_n358_n500# w_n394_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__nfet_01v8_AH5E2K a_500_n500# a_n558_n500# a_n500_n588# VSUBS
X0 a_500_n500# a_n500_n588# a_n558_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__nfet_01v8_QP5WRD a_500_n2936# a_500_n5372# a_n500_n1806# a_500_718#
+ a_n500_3066# a_n500_n4242# a_n500_630# a_n500_n6678# a_n558_1936# a_n558_4372# a_n558_n9026#
+ a_n558_n6590# a_500_n500# a_500_6808# a_n500_6720# a_500_3154# a_500_n7808# a_n500_n9114#
+ a_500_n4154# a_500_n1718# a_n558_n500# a_n500_n3024# a_n558_6808# a_n558_n2936#
+ a_n558_3154# a_n558_n5372# a_n558_718# a_n500_n588# a_n500_5502# a_500_8026# a_500_5590#
+ a_n500_7938# a_500_n9026# a_n500_1848# a_500_n6590# a_n500_4284# a_n500_n5460# a_n558_n7808#
+ a_n500_n7896# a_n558_8026# a_n558_n1718# a_n558_5590# a_n558_n4154# a_500_1936#
+ a_500_4372# VSUBS
X0 a_500_4372# a_n500_4284# a_n558_4372# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1 a_500_n6590# a_n500_n6678# a_n558_n6590# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X2 a_500_5590# a_n500_5502# a_n558_5590# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X3 a_500_n1718# a_n500_n1806# a_n558_n1718# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X4 a_500_n2936# a_n500_n3024# a_n558_n2936# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X5 a_500_n4154# a_n500_n4242# a_n558_n4154# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X6 a_500_718# a_n500_630# a_n558_718# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X7 a_500_n5372# a_n500_n5460# a_n558_n5372# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X8 a_500_6808# a_n500_6720# a_n558_6808# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X9 a_500_8026# a_n500_7938# a_n558_8026# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X10 a_500_n500# a_n500_n588# a_n558_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X11 a_500_1936# a_n500_1848# a_n558_1936# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X12 a_500_n7808# a_n500_n7896# a_n558_n7808# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X13 a_500_3154# a_n500_3066# a_n558_3154# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X14 a_500_n9026# a_n500_n9114# a_n558_n9026# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__pfet_01v8_UDM5A5 a_n558_n7916# a_n500_5583# a_500_1972# a_n558_8152#
+ a_n500_8055# a_500_4444# w_n594_3108# w_n594_6816# a_500_n2972# a_500_736# a_500_n5444#
+ a_n500_n597# w_n594_636# a_500_n500# w_n594_n3072# a_n558_1972# w_n594_n6780# w_n594_n600#
+ a_n500_1875# a_n558_4444# w_n594_n9252# a_n500_4347# a_n558_n6680# a_n558_n9152#
+ a_n500_n5541# a_n500_639# a_500_3208# a_n500_n8013# a_500_6916# a_500_n1736# a_n558_n500#
+ a_500_n4208# w_n594_5580# a_500_n7916# w_n594_8052# w_n594_n5544# a_n558_736# a_n558_3208#
+ w_n594_n8016# a_n558_n2972# a_n558_6916# a_n558_n5444# a_n500_n1833# a_n500_6819#
+ a_n500_n4305# w_n594_1872# a_500_5680# a_n500_n3069# w_n594_4344# a_n500_n6777#
+ a_500_8152# w_n594_n1836# a_n500_n9249# a_500_n6680# w_n594_n4308# a_n500_3111#
+ a_500_n9152# a_n558_n1736# a_n558_n4208# a_n558_5680#
X0 a_500_1972# a_n500_1875# a_n558_1972# w_n594_1872# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1 a_500_6916# a_n500_6819# a_n558_6916# w_n594_6816# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X2 a_500_4444# a_n500_4347# a_n558_4444# w_n594_4344# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X3 a_500_n9152# a_n500_n9249# a_n558_n9152# w_n594_n9252# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X4 a_500_3208# a_n500_3111# a_n558_3208# w_n594_3108# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X5 a_500_n2972# a_n500_n3069# a_n558_n2972# w_n594_n3072# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X6 a_500_n7916# a_n500_n8013# a_n558_n7916# w_n594_n8016# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X7 a_500_n5444# a_n500_n5541# a_n558_n5444# w_n594_n5544# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X8 a_500_n500# a_n500_n597# a_n558_n500# w_n594_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X9 a_500_n1736# a_n500_n1833# a_n558_n1736# w_n594_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X10 a_500_n4208# a_n500_n4305# a_n558_n4208# w_n594_n4308# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X11 a_500_736# a_n500_639# a_n558_736# w_n594_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X12 a_500_n6680# a_n500_n6777# a_n558_n6680# w_n594_n6780# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X13 a_500_5680# a_n500_5583# a_n558_5680# w_n594_5580# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X14 a_500_8152# a_n500_8055# a_n558_8152# w_n594_8052# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__nfet_01v8_3ZAA45 a_100_n500# a_n158_n500# a_n100_n588# VSUBS
X0 a_100_n500# a_n100_n588# a_n158_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=1
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__pfet_01v8_SKU9VM a_n500_n597# a_500_n500# w_n594_n600# a_n558_n500#
X0 a_500_n500# a_n500_n597# a_n558_n500# w_n594_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__pfet_01v8_E769TZ a_n1558_11242# a_n1558_n14714# a_n1500_n43239#
+ w_n1594_n3690# a_n1500_n11103# a_n1558_50794# a_1500_n23366# a_n1500_n50655# w_n1594_n56838#
+ w_n1594_n24702# a_1500_n30782# a_n1500_3729# a_n1558_n60446# w_n1594_12378# w_n1594_n63018#
+ a_1500_n8534# a_n1558_14950# a_1500_n19658# a_n1500_n14811# a_n1500_n46947# w_n1594_9906#
+ w_n1594_n6162# a_1500_22366# a_n1500_22269# a_n1558_53266# a_n1558_n56738# a_n1558_n24602#
+ a_n1558_21130# a_n1500_n53127# w_n1594_n13578# a_n1558_60682# a_1500_n33254# a_n1500_n60543#
+ w_n1594_n20994# a_1500_n40670# a_1500_18658# a_n1558_49558# a_n1558_17422# w_n1594_22266#
+ a_n1500_n49419# w_n1594_n9870# a_n1500_25977# a_n1558_56974# a_n1500_n56835# a_1500_n29546#
+ a_n1558_n3590# a_1500_n36962# a_n1500_9909# a_n1558_n13478# a_1500_32254# a_n1500_32157#
+ a_n1558_n20894# a_n1500_n63015# w_n1594_18558# w_n1594_n23466# a_1500_n43142# w_n1594_n30882#
+ w_n1594_25974# a_n1500_n2451# a_1500_28546# a_1500_n7298# a_n1500_28449# a_n1558_59446#
+ a_n1558_27310# a_n1500_n13575# a_n1500_n59307# w_n1594_32154# w_n1594_n19758# a_1500_35962#
+ a_n1558_n6062# a_n1500_35865# a_1500_n39434# a_n1500_n20991# a_n1558_n23366# a_1500_n46850#
+ a_1500_42142# a_n1500_42045# a_n1558_n30782# w_n1594_n33354# w_n1594_28446# a_1500_n53030#
+ w_n1594_n40770# w_n1594_35862# a_n1558_n9770# w_n1594_18# a_n1558_16186# a_n1500_21#
+ a_n1558_n19658# a_n1500_n16047# a_1500_38434# a_n1500_38337# a_n1500_n55599# a_n1500_n23463#
+ w_n1594_n29646# a_1500_45850# w_n1594_42042# a_n1500_45753# a_n1558_40906# a_1500_n49322#
+ a_n1558_n33254# a_1500_52030# a_n1500_n8631# a_n1558_n40670# a_n1558_19894# w_n1594_n43242#
+ a_n1500_n19755# w_n1594_38334# w_n1594_45750# a_n1558_26074# a_n1558_n29546# a_1500_48322#
+ a_n1500_48225# a_1500_n38198# a_n1558_33490# a_n1558_n36962# a_n1500_n33351# w_n1594_n39534#
+ a_n1500_55641# a_1500_n59210# w_n1594_n46950# a_1500_n62918# a_n1558_n43142# a_n1558_29782#
+ w_n1594_n53130# a_n1500_n29643# w_n1594_48222# a_1500_37198# a_n1558_n39434# a_1500_58210#
+ a_n1500_58113# a_n1500_12381# a_1500_n1118# a_1500_n48086# a_n1558_n46850# a_1500_61918#
+ w_n1594_n49422# a_n1500_n7395# a_n1558_n53030# w_n1594_37098# a_n1558_39670# a_n1500_n39531#
+ w_n1594_58110# a_1500_n4826# w_n1594_61818# a_1500_47086# a_n1558_10006# a_n1558_n49322#
+ w_n1594_n2454# w_n1594_n38298# a_1500_2590# w_n1594_2490# w_n1594_n59310# a_n1500_6201#
+ a_n1500_18561# a_n1558_13714# a_n1558_2590# a_1500_n25838# a_n1558_n38198# a_1500_5062#
+ a_1500_118# a_n1558_n59210# w_n1594_n48186# w_n1594_n16050# a_n1558_n62918# a_1500_n32018#
+ a_n1500_2493# a_1500_24838# a_n1558_5062# a_n1500_n38295# w_n1594_n8634# a_1500_8770#
+ a_n1558_55738# a_n1558_23602# a_n1558_n2354# w_n1594_8670# a_1500_n35726# a_n1558_n48086#
+ a_1500_31018# w_n1594_n58074# w_n1594_24738# a_n1558_8770# a_n1500_n1215# a_n1558_12478#
+ a_n1500_n12339# a_n1500_n48183# a_1500_34726# a_n1500_34629# w_n1594_n25938# a_1500_n45614#
+ a_n1500_8673# w_n1594_n32118# a_n1500_n4923# w_n1594_34626# a_n1558_n8534# w_n1594_n7398#
+ a_n1558_22366# a_n1558_n25838# a_n1500_n22227# a_n1500_n58071# a_1500_44614# a_n1500_44517#
+ a_n1500_n61779# w_n1594_n35826# a_n1500_51933# a_1500_n55502# a_n1558_n32018# a_n1558_18658#
+ w_n1594_n42006# a_n1500_n18519# a_n1500_n25935# w_n1594_44514# w_n1594_51930# a_n1558_32254#
+ a_n1558_n35726# a_n1500_n32115# a_1500_54502# a_n1500_54405# a_1500_n44378# a_1500_n12242#
+ w_n1594_n45714# a_n1500_61821# a_1500_n51794# a_n1500_n3687# a_n1558_28546# a_n1558_n7298#
+ a_n1500_n28407# a_n1558_35962# a_n1500_n35823# w_n1594_54402# a_1500_n15950# a_1500_43378#
+ a_1500_11242# a_n1500_11145# a_n1558_42142# a_n1558_n45614# a_1500_50794# a_n1500_n42003#
+ a_n1500_50697# a_1500_n54266# a_1500_n22130# a_n1500_n6159# w_n1594_n55602# a_1500_n61682#
+ a_n1558_38434# a_n1500_n24699# w_n1594_43278# w_n1594_11142# a_1500_14950# a_n1500_46989#
+ a_n1558_45850# a_n1500_14853# a_1500_n18422# a_n1500_n45711# w_n1594_50694# a_1500_n57974#
+ a_n1500_n9867# w_n1594_n1218# a_1500_53266# a_1500_1354# a_n1500_53169# a_1500_21130#
+ a_n1500_21033# a_n1558_n55502# a_n1558_52030# w_n1594_1254# w_n1594_n12342# w_n1594_n44478#
+ a_1500_60682# a_n1500_60585# w_n1594_14850# w_n1594_n51894# w_n1594_46986# a_1500_49558#
+ a_1500_17422# a_n1558_48322# a_n1500_17325# a_n1500_n34587# a_1500_56974# a_n1558_1354#
+ w_n1594_53166# w_n1594_21030# w_n1594_n4926# a_n1500_56877# a_n1500_24741# a_1500_n3590#
+ a_1500_n28310# w_n1594_60582# w_n1594_4962# a_n1558_n44378# a_n1558_n12242# a_n1558_n51794#
+ w_n1594_17322# w_n1594_n22230# w_n1594_n54366# w_n1594_49458# a_n1500_1257# w_n1594_n61782#
+ w_n1594_56874# a_n1558_37198# a_n1500_n37059# a_1500_59446# a_1500_27310# a_1500_7534#
+ a_n1500_59349# a_n1500_27213# a_1500_n6062# a_1500_n17186# a_n1558_58210# a_n1558_n15950#
+ a_n1500_n44475# a_n1558_n1118# w_n1594_7434# w_n1594_n18522# a_n1558_61918# a_n1500_n51891#
+ a_n1558_n54266# a_1500_n41906# a_n1500_4965# a_n1558_n22130# a_n1558_n61682# w_n1594_59346#
+ w_n1594_27210# a_n1558_7534# a_1500_n9770# w_n1594_30918# a_n1558_n4826# a_1500_16186#
+ a_n1500_16089# a_n1558_47086# a_n1558_n18422# a_n1500_37101# a_n1558_n57974# a_1500_n27074#
+ a_n1500_n54363# a_1500_40906# w_n1594_n28410# a_n1500_40809# a_1500_n34490# a_n1500_7437#
+ w_n1594_16086# a_1500_19894# a_n1500_19797# w_n1594_40806# a_1500_26074# a_1500_6298#
+ a_n1558_n28310# w_n1594_6198# w_n1594_n17286# a_1500_33490# a_n1500_33393# w_n1594_19794#
+ a_n1558_6298# a_1500_29782# a_n1500_29685# a_n1558_24838# w_n1594_33390# a_n1558_n17186#
+ a_n1558_118# a_n1558_31018# w_n1594_n27174# a_n1500_43281# a_n1558_n41906# a_1500_n11006#
+ w_n1594_29682# w_n1594_n34590# a_1500_n50558# a_n1500_n17283# a_1500_39670# a_n1500_39573#
+ a_n1558_34726# a_1500_n14714# a_n1558_n27074# a_1500_10006# a_n1558_n34490# w_n1594_n37062#
+ w_n1594_39570# a_1500_n60446# a_n1500_n27171# a_1500_13714# a_n1500_13617# a_n1500_49461#
+ a_n1558_44614# a_n1500_n30879# a_1500_n56738# a_1500_n24602# w_n1594_n11106# w_n1594_n50658#
+ w_n1594_13614# a_1500_55738# a_1500_23602# a_1500_3826# a_n1500_23505# a_1500_n2354#
+ a_1500_n13478# a_n1558_54502# a_n1500_n40767# w_n1594_3726# w_n1594_n14814# a_n1500_30921#
+ a_1500_n20894# a_n1558_n11006# a_n1558_n50558# w_n1594_n60546# a_n1558_3826# w_n1594_55638#
+ w_n1594_23502# a_1500_12478# a_n1558_43378#
X0 a_1500_53266# a_n1500_53169# a_n1558_53266# w_n1594_53166# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1 a_1500_n18422# a_n1500_n18519# a_n1558_n18422# w_n1594_n18522# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X2 a_1500_n45614# a_n1500_n45711# a_n1558_n45614# w_n1594_n45714# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X3 a_1500_n43142# a_n1500_n43239# a_n1558_n43142# w_n1594_n43242# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X4 a_1500_n22130# a_n1500_n22227# a_n1558_n22130# w_n1594_n22230# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X5 a_1500_n3590# a_n1500_n3687# a_n1558_n3590# w_n1594_n3690# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X6 a_1500_35962# a_n1500_35865# a_n1558_35962# w_n1594_35862# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X7 a_1500_33490# a_n1500_33393# a_n1558_33490# w_n1594_33390# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X8 a_1500_60682# a_n1500_60585# a_n1558_60682# w_n1594_60582# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X9 a_1500_12478# a_n1500_12381# a_n1558_12478# w_n1594_12378# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X10 a_1500_38434# a_n1500_38337# a_n1558_38434# w_n1594_38334# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X11 a_1500_6298# a_n1500_6201# a_n1558_6298# w_n1594_6198# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X12 a_1500_n55502# a_n1500_n55599# a_n1558_n55502# w_n1594_n55602# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X13 a_1500_n32018# a_n1500_n32115# a_n1558_n32018# w_n1594_n32118# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X14 a_1500_45850# a_n1500_45753# a_n1558_45850# w_n1594_45750# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X15 a_1500_24838# a_n1500_24741# a_n1558_24838# w_n1594_24738# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X16 a_1500_n38198# a_n1500_n38295# a_n1558_n38198# w_n1594_n38298# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X17 a_1500_22366# a_n1500_22269# a_n1558_22366# w_n1594_22266# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X18 a_1500_48322# a_n1500_48225# a_n1558_48322# w_n1594_48222# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X19 a_1500_n14714# a_n1500_n14811# a_n1558_n14714# w_n1594_n14814# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X20 a_1500_n41906# a_n1500_n42003# a_n1558_n41906# w_n1594_n42006# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X21 a_1500_n12242# a_n1500_n12339# a_n1558_n12242# w_n1594_n12342# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X22 a_1500_34726# a_n1500_34629# a_n1558_34726# w_n1594_34626# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X23 a_1500_61918# a_n1500_61821# a_n1558_61918# w_n1594_61818# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X24 a_1500_32254# a_n1500_32157# a_n1558_32254# w_n1594_32154# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X25 a_1500_n48086# a_n1500_n48183# a_n1558_n48086# w_n1594_n48186# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X26 a_1500_58210# a_n1500_58113# a_n1558_58210# w_n1594_58110# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X27 a_1500_n24602# a_n1500_n24699# a_n1558_n24602# w_n1594_n24702# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X28 a_1500_14950# a_n1500_14853# a_n1558_14950# w_n1594_14850# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X29 a_1500_n8534# a_n1500_n8631# a_n1558_n8534# w_n1594_n8634# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X30 a_1500_n57974# a_n1500_n58071# a_n1558_n57974# w_n1594_n58074# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X31 a_1500_n6062# a_n1500_n6159# a_n1558_n6062# w_n1594_n6162# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X32 a_1500_n34490# a_n1500_n34587# a_n1558_n34490# w_n1594_n34590# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X33 a_1500_17422# a_n1500_17325# a_n1558_17422# w_n1594_17322# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X34 a_1500_44614# a_n1500_44517# a_n1558_44614# w_n1594_44514# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X35 a_1500_42142# a_n1500_42045# a_n1558_42142# w_n1594_42042# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X36 a_1500_8770# a_n1500_8673# a_n1558_8770# w_n1594_8670# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X37 a_1500_n11006# a_n1500_n11103# a_n1558_n11006# w_n1594_n11106# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X38 a_1500_n19658# a_n1500_n19755# a_n1558_n19658# w_n1594_n19758# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X39 a_1500_n46850# a_n1500_n46947# a_n1558_n46850# w_n1594_n46950# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X40 a_1500_n17186# a_n1500_n17283# a_n1558_n17186# w_n1594_n17286# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X41 a_1500_27310# a_n1500_27213# a_n1558_27310# w_n1594_27210# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X42 a_1500_n44378# a_n1500_n44475# a_n1558_n44378# w_n1594_n44478# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X43 a_1500_54502# a_n1500_54405# a_n1558_54502# w_n1594_54402# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X44 a_1500_52030# a_n1500_51933# a_n1558_52030# w_n1594_51930# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X45 a_1500_31018# a_n1500_30921# a_n1558_31018# w_n1594_30918# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X46 a_1500_n4826# a_n1500_n4923# a_n1558_n4826# w_n1594_n4926# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X47 a_1500_37198# a_n1500_37101# a_n1558_37198# w_n1594_37098# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X48 a_1500_n2354# a_n1500_n2451# a_n1558_n2354# w_n1594_n2454# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X49 a_1500_n51794# a_n1500_n51891# a_n1558_n51794# w_n1594_n51894# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X50 a_1500_n29546# a_n1500_n29643# a_n1558_n29546# w_n1594_n29646# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X51 a_1500_13714# a_n1500_13617# a_n1558_13714# w_n1594_13614# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X52 a_1500_n56738# a_n1500_n56835# a_n1558_n56738# w_n1594_n56838# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X53 a_1500_11242# a_n1500_11145# a_n1558_11242# w_n1594_11142# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X54 a_1500_40906# a_n1500_40809# a_n1558_40906# w_n1594_40806# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X55 a_1500_n27074# a_n1500_n27171# a_n1558_n27074# w_n1594_n27174# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X56 a_1500_n54266# a_n1500_n54363# a_n1558_n54266# w_n1594_n54366# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X57 a_1500_19894# a_n1500_19797# a_n1558_19894# w_n1594_19794# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X58 a_1500_2590# a_n1500_2493# a_n1558_2590# w_n1594_2490# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X59 a_1500_n59210# a_n1500_n59307# a_n1558_n59210# w_n1594_n59310# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X60 a_1500_7534# a_n1500_7437# a_n1558_7534# w_n1594_7434# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X61 a_1500_49558# a_n1500_49461# a_n1558_49558# w_n1594_49458# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X62 a_1500_n36962# a_n1500_n37059# a_n1558_n36962# w_n1594_n37062# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X63 a_1500_5062# a_n1500_4965# a_n1558_5062# w_n1594_4962# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X64 a_1500_47086# a_n1500_46989# a_n1558_47086# w_n1594_46986# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X65 a_1500_n15950# a_n1500_n16047# a_n1558_n15950# w_n1594_n16050# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X66 a_1500_n61682# a_n1500_n61779# a_n1558_n61682# w_n1594_n61782# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X67 a_1500_n13478# a_n1500_n13575# a_n1558_n13478# w_n1594_n13578# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X68 a_1500_23602# a_n1500_23505# a_n1558_23602# w_n1594_23502# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X69 a_1500_n40670# a_n1500_n40767# a_n1558_n40670# w_n1594_n40770# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X70 a_1500_n39434# a_n1500_n39531# a_n1558_n39434# w_n1594_n39534# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X71 a_1500_21130# a_n1500_21033# a_n1558_21130# w_n1594_21030# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X72 a_1500_29782# a_n1500_29685# a_n1558_29782# w_n1594_29682# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X73 a_1500_56974# a_n1500_56877# a_n1558_56974# w_n1594_56874# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X74 a_1500_59446# a_n1500_59349# a_n1558_59446# w_n1594_59346# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X75 a_1500_n20894# a_n1500_n20991# a_n1558_n20894# w_n1594_n20994# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X76 a_1500_n25838# a_n1500_n25935# a_n1558_n25838# w_n1594_n25938# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X77 a_1500_n23366# a_n1500_n23463# a_n1558_n23366# w_n1594_n23466# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X78 a_1500_n50558# a_n1500_n50655# a_n1558_n50558# w_n1594_n50658# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X79 a_1500_n49322# a_n1500_n49419# a_n1558_n49322# w_n1594_n49422# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X80 a_1500_n1118# a_n1500_n1215# a_n1558_n1118# w_n1594_n1218# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X81 a_1500_n9770# a_n1500_n9867# a_n1558_n9770# w_n1594_n9870# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X82 a_1500_n28310# a_n1500_n28407# a_n1558_n28310# w_n1594_n28410# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X83 a_1500_n7298# a_n1500_n7395# a_n1558_n7298# w_n1594_n7398# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X84 a_1500_10006# a_n1500_9909# a_n1558_10006# w_n1594_9906# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X85 a_1500_39670# a_n1500_39573# a_n1558_39670# w_n1594_39570# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X86 a_1500_18658# a_n1500_18561# a_n1558_18658# w_n1594_18558# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X87 a_1500_n53030# a_n1500_n53127# a_n1558_n53030# w_n1594_n53130# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X88 a_1500_3826# a_n1500_3729# a_n1558_3826# w_n1594_3726# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X89 a_1500_16186# a_n1500_16089# a_n1558_16186# w_n1594_16086# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X90 a_1500_1354# a_n1500_1257# a_n1558_1354# w_n1594_1254# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X91 a_1500_43378# a_n1500_43281# a_n1558_43378# w_n1594_43278# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X92 a_1500_n30782# a_n1500_n30879# a_n1558_n30782# w_n1594_n30882# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X93 a_1500_118# a_n1500_21# a_n1558_118# w_n1594_18# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X94 a_1500_n35726# a_n1500_n35823# a_n1558_n35726# w_n1594_n35826# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X95 a_1500_n62918# a_n1500_n63015# a_n1558_n62918# w_n1594_n63018# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X96 a_1500_n33254# a_n1500_n33351# a_n1558_n33254# w_n1594_n33354# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X97 a_1500_n60446# a_n1500_n60543# a_n1558_n60446# w_n1594_n60546# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X98 a_1500_50794# a_n1500_50697# a_n1558_50794# w_n1594_50694# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X99 a_1500_28546# a_n1500_28449# a_n1558_28546# w_n1594_28446# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X100 a_1500_55738# a_n1500_55641# a_n1558_55738# w_n1594_55638# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X101 a_1500_26074# a_n1500_25977# a_n1558_26074# w_n1594_25974# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__pfet_01v8_UDMRD5 a_n558_n10388# a_n558_n7916# a_n500_5583# a_n500_n10485#
+ a_500_1972# a_n558_8152# a_n500_8055# a_500_4444# w_n594_3108# w_n594_6816# a_500_n2972#
+ a_500_736# a_500_n5444# a_n500_n597# w_n594_636# a_500_n500# a_500_9388# w_n594_n3072#
+ a_n558_1972# w_n594_n6780# w_n594_n600# a_n500_1875# a_n558_4444# w_n594_n9252#
+ a_n500_4347# a_n558_n6680# w_n594_n10488# a_n558_n9152# a_n500_n5541# a_n500_639#
+ a_500_3208# a_n500_n8013# a_500_6916# a_500_n1736# a_n558_n500# a_n558_9388# a_500_n4208#
+ w_n594_5580# a_500_n7916# w_n594_8052# w_n594_n5544# a_n558_736# a_n558_3208# w_n594_n8016#
+ a_n558_n2972# a_n558_6916# a_n558_n5444# a_n500_n1833# a_n500_6819# a_n500_n4305#
+ w_n594_1872# a_500_5680# a_n500_9291# a_n500_n3069# w_n594_4344# a_n500_n6777# a_500_8152#
+ w_n594_n1836# a_n500_n9249# a_500_n6680# w_n594_n4308# a_500_n10388# a_n500_3111#
+ a_500_n9152# a_n558_n1736# w_n594_9288# a_n558_n4208# a_n558_5680#
X0 a_500_1972# a_n500_1875# a_n558_1972# w_n594_1872# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1 a_500_6916# a_n500_6819# a_n558_6916# w_n594_6816# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X2 a_500_4444# a_n500_4347# a_n558_4444# w_n594_4344# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X3 a_500_n9152# a_n500_n9249# a_n558_n9152# w_n594_n9252# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X4 a_500_3208# a_n500_3111# a_n558_3208# w_n594_3108# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X5 a_500_n2972# a_n500_n3069# a_n558_n2972# w_n594_n3072# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X6 a_500_n7916# a_n500_n8013# a_n558_n7916# w_n594_n8016# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X7 a_500_9388# a_n500_9291# a_n558_9388# w_n594_9288# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X8 a_500_n5444# a_n500_n5541# a_n558_n5444# w_n594_n5544# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X9 a_500_n500# a_n500_n597# a_n558_n500# w_n594_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X10 a_500_n1736# a_n500_n1833# a_n558_n1736# w_n594_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X11 a_500_n4208# a_n500_n4305# a_n558_n4208# w_n594_n4308# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X12 a_500_n10388# a_n500_n10485# a_n558_n10388# w_n594_n10488# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X13 a_500_736# a_n500_639# a_n558_736# w_n594_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X14 a_500_n6680# a_n500_n6777# a_n558_n6680# w_n594_n6780# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X15 a_500_5680# a_n500_5583# a_n558_5680# w_n594_5580# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X16 a_500_8152# a_n500_8055# a_n558_8152# w_n594_8052# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__pfet_01v8_RRU5GE a_n300_n1833# w_n394_n1836# a_n358_n1736# a_300_736#
+ w_n394_636# a_n300_n597# a_300_n500# a_n300_639# w_n394_n600# a_300_n1736# a_n358_n500#
+ a_n358_736#
X0 a_300_n500# a_n300_n597# a_n358_n500# w_n394_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X1 a_300_736# a_n300_639# a_n358_736# w_n394_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X2 a_300_n1736# a_n300_n1833# a_n358_n1736# w_n394_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__pfet_01v8_SLZ774 w_n1594_n600# a_n1500_n597# a_1500_n500# a_n1558_n500#
X0 a_1500_n500# a_n1500_n597# a_n1558_n500# w_n1594_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
.ends

.subckt opamp_cascode IN_P IN_M VCC VSS OUT VB_A VB_B IB
Xsky130_fd_pr__nfet_01v8_SCE452_3 VSS bias21 bias21 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM9_dummy_15 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM5_1 VCC IN_M IN_M bias3 VCC VCC m1_44990_37960# m1_44990_37960# m1_44990_37960#
+ bias3 IN_M bias3 m1_44990_37960# bias3 IN_M m1_44990_37960# bias3 VCC IN_M IN_M
+ bias3 VCC IN_M IN_M IN_M VCC VCC VCC IN_M IN_M IN_M m1_44990_37960# m1_44990_37960#
+ m1_44990_37960# bias3 IN_M VCC bias3 m1_44990_37960# bias3 m1_44990_37960# IN_M
+ VCC bias3 m1_44990_37960# VCC bias3 VCC VCC m1_44990_37960# bias3 m1_44990_37960#
+ bias3 bias3 m1_44990_37960# bias3 VCC m1_44990_37960# IN_M VCC sky130_fd_pr__pfet_01v8_7DHACV
XXM4_dummy_2 dummy_4 bias3 dummy_4 dummy_4 bias3 dummy_4 bias3 dummy_4 bias3 dummy_4
+ dummy_4 dummy_4 dummy_4 dummy_4 bias3 dummy_4 dummy_4 bias3 VSS sky130_fd_pr__nfet_01v8_MHE452
XXM9_dummy_16 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM100_4 IB VCC IB IB VCC VCC VCC IB sky130_fd_pr__pfet_01v8_P2UXFR
XXM4_dummy_3 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM9_dummy_17 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_dummy_18 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
Xsky130_fd_pr__nfet_01v8_VT3ZQW_0 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM9_dummy_19 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
Xsky130_fd_pr__pfet_01v8_RRUZAE_0 dummy_100 IB IB VCC VCC dummy_100 dummy_100 dummy_100
+ dummy_100 VCC VCC IB dummy_100 IB dummy_100 IB VCC dummy_100 dummy_100 dummy_100
+ sky130_fd_pr__pfet_01v8_RRUZAE
XXM4_dummy_7 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
Xsky130_fd_pr__pfet_01v8_P2UXFR_0 IB VCC VCC IB IB VCC IB VCC sky130_fd_pr__pfet_01v8_P2UXFR
Xsky130_fd_pr__pfet_01v8_ZLZ7XS_0 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM100_dummy_1 dummy_100 IB IB VCC VCC dummy_100 dummy_100 dummy_100 dummy_100 VCC
+ VCC IB dummy_100 IB dummy_100 IB VCC dummy_100 dummy_100 dummy_100 sky130_fd_pr__pfet_01v8_RRUZAE
XXM1_1 m1m2 m1m2 bias1 VCC bias1 m1m2 VCC bias1 VCC VCC VCC bias1 m1m2 VCC VCC m1m2
+ VCC bias1 bias1 VCC VCC VCC bias1 m1m2 m1m2 m1m2 m1m2 bias1 VCC m1m2 VCC bias1 VCC
+ VCC VCC m1m2 m1m2 VCC bias1 VCC bias1 m1m2 bias1 VCC m1m2 VCC bias1 m1m2 VCC bias1
+ m1m2 VCC VCC VCC VCC VCC bias1 VCC VCC bias1 m1m2 m1m2 bias1 bias1 VCC VCC VCC m1m2
+ bias1 VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC VCC VCC VCC VCC m1m2 VCC m1m2 bias1
+ m1m2 bias1 VCC bias1 bias1 bias1 VCC VCC VCC bias1 m1m2 VCC m1m2 VCC bias1 m1m2
+ m1m2 VCC VCC bias1 VCC m1m2 m1m2 VCC bias1 VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC
+ m1m2 m1m2 VCC bias1 VCC VCC m1m2 VCC bias1 bias1 VCC VCC m1m2 VCC bias1 m1m2 VCC
+ m1m2 bias1 VCC VCC VCC m1m2 m1m2 VCC VCC VCC VCC VCC bias1 bias1 m1m2 m1m2 VCC m1m2
+ VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 bias1 VCC VCC m1m2 m1m2 m1m2 VCC VCC m1m2
+ VCC VCC VCC m1m2 bias1 m1m2 bias1 bias1 VCC bias1 VCC VCC bias1 VCC bias1 VCC m1m2
+ VCC m1m2 m1m2 bias1 bias1 VCC bias1 bias1 VCC bias1 VCC m1m2 m1m2 VCC bias1 bias1
+ VCC VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC VCC VCC bias1 m1m2 m1m2 bias1 m1m2 bias1
+ VCC VCC VCC VCC bias1 m1m2 m1m2 VCC bias1 bias1 VCC VCC bias1 VCC VCC m1m2 bias1
+ VCC VCC VCC bias1 m1m2 bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC bias1 VCC bias1
+ m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC VCC VCC VCC m1m2 bias1 bias1 VCC m1m2 VCC
+ VCC VCC bias1 bias1 VCC VCC VCC VCC m1m2 m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC
+ m1m2 bias1 VCC VCC VCC bias1 bias1 VCC VCC m1m2 m1m2 bias1 m1m2 VCC VCC bias1 m1m2
+ VCC bias1 m1m2 m1m2 VCC VCC m1m2 VCC VCC m1m2 VCC bias1 m1m2 m1m2 bias1 m1m2 VCC
+ bias1 VCC VCC bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC m1m2 VCC VCC VCC bias1 VCC
+ m1m2 VCC bias1 m1m2 VCC m1m2 m1m2 m1m2 VCC bias1 m1m2 VCC VCC VCC VCC bias1 VCC
+ bias1 m1m2 VCC m1m2 VCC m1m2 VCC VCC VCC bias1 VCC bias1 bias1 m1m2 bias1 VCC VCC
+ VCC VCC VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC bias1 VCC m1m2 m1m2 VCC
+ m1m2 VCC VCC VCC m1m2 sky130_fd_pr__pfet_01v8_F76D73
XXM4_dummy_9 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM1_2 m1m2 m1m2 bias1 VCC bias1 m1m2 VCC bias1 VCC VCC VCC bias1 m1m2 VCC VCC m1m2
+ VCC bias1 bias1 VCC VCC VCC bias1 m1m2 m1m2 m1m2 m1m2 bias1 VCC m1m2 VCC bias1 VCC
+ VCC VCC m1m2 m1m2 VCC bias1 VCC bias1 m1m2 bias1 VCC m1m2 VCC bias1 m1m2 VCC bias1
+ m1m2 VCC VCC VCC VCC VCC bias1 VCC VCC bias1 m1m2 m1m2 bias1 bias1 VCC VCC VCC m1m2
+ bias1 VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC VCC VCC VCC VCC m1m2 VCC m1m2 bias1
+ m1m2 bias1 VCC bias1 bias1 bias1 VCC VCC VCC bias1 m1m2 VCC m1m2 VCC bias1 m1m2
+ m1m2 VCC VCC bias1 VCC m1m2 m1m2 VCC bias1 VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC
+ m1m2 m1m2 VCC bias1 VCC VCC m1m2 VCC bias1 bias1 VCC VCC m1m2 VCC bias1 m1m2 VCC
+ m1m2 bias1 VCC VCC VCC m1m2 m1m2 VCC VCC VCC VCC VCC bias1 bias1 m1m2 m1m2 VCC m1m2
+ VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 bias1 VCC VCC m1m2 m1m2 m1m2 VCC VCC m1m2
+ VCC VCC VCC m1m2 bias1 m1m2 bias1 bias1 VCC bias1 VCC VCC bias1 VCC bias1 VCC m1m2
+ VCC m1m2 m1m2 bias1 bias1 VCC bias1 bias1 VCC bias1 VCC m1m2 m1m2 VCC bias1 bias1
+ VCC VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC VCC VCC bias1 m1m2 m1m2 bias1 m1m2 bias1
+ VCC VCC VCC VCC bias1 m1m2 m1m2 VCC bias1 bias1 VCC VCC bias1 VCC VCC m1m2 bias1
+ VCC VCC VCC bias1 m1m2 bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC bias1 VCC bias1
+ m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC VCC VCC VCC m1m2 bias1 bias1 VCC m1m2 VCC
+ VCC VCC bias1 bias1 VCC VCC VCC VCC m1m2 m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC
+ m1m2 bias1 VCC VCC VCC bias1 bias1 VCC VCC m1m2 m1m2 bias1 m1m2 VCC VCC bias1 m1m2
+ VCC bias1 m1m2 m1m2 VCC VCC m1m2 VCC VCC m1m2 VCC bias1 m1m2 m1m2 bias1 m1m2 VCC
+ bias1 VCC VCC bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC m1m2 VCC VCC VCC bias1 VCC
+ m1m2 VCC bias1 m1m2 VCC m1m2 m1m2 m1m2 VCC bias1 m1m2 VCC VCC VCC VCC bias1 VCC
+ bias1 m1m2 VCC m1m2 VCC m1m2 VCC VCC VCC bias1 VCC bias1 bias1 m1m2 bias1 VCC VCC
+ VCC VCC VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC bias1 VCC m1m2 m1m2 VCC
+ m1m2 VCC VCC VCC m1m2 sky130_fd_pr__pfet_01v8_F76D73
XXM100_dummy_3 IB VCC dummy_100 IB dummy_100 VCC dummy_100 dummy_100 sky130_fd_pr__pfet_01v8_P2UXFR
XXM3_dummy_1 VB_B dummy_3 dummy_3 dummy_3 VB_B dummy_3 VB_B VB_B VB_B VB_B dummy_3
+ dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 VB_B dummy_3 dummy_3 dummy_3 VB_B dummy_3
+ dummy_3 dummy_3 VB_B dummy_3 dummy_3 dummy_3 dummy_3 VB_B dummy_3 dummy_3 VB_B VB_B
+ dummy_3 dummy_3 VB_B dummy_3 VB_B dummy_3 VB_B VB_B dummy_3 VB_B dummy_3 dummy_3
+ dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 VSS sky130_fd_pr__nfet_01v8_WK8VRD
XXM1_3 m1m2 m1m2 bias1 VCC bias1 m1m2 VCC bias1 VCC VCC VCC bias1 m1m2 VCC VCC m1m2
+ VCC bias1 bias1 VCC VCC VCC bias1 m1m2 m1m2 m1m2 m1m2 bias1 VCC m1m2 VCC bias1 VCC
+ VCC VCC m1m2 m1m2 VCC bias1 VCC bias1 m1m2 bias1 VCC m1m2 VCC bias1 m1m2 VCC bias1
+ m1m2 VCC VCC VCC VCC VCC bias1 VCC VCC bias1 m1m2 m1m2 bias1 bias1 VCC VCC VCC m1m2
+ bias1 VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC VCC VCC VCC VCC m1m2 VCC m1m2 bias1
+ m1m2 bias1 VCC bias1 bias1 bias1 VCC VCC VCC bias1 m1m2 VCC m1m2 VCC bias1 m1m2
+ m1m2 VCC VCC bias1 VCC m1m2 m1m2 VCC bias1 VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC
+ m1m2 m1m2 VCC bias1 VCC VCC m1m2 VCC bias1 bias1 VCC VCC m1m2 VCC bias1 m1m2 VCC
+ m1m2 bias1 VCC VCC VCC m1m2 m1m2 VCC VCC VCC VCC VCC bias1 bias1 m1m2 m1m2 VCC m1m2
+ VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 bias1 VCC VCC m1m2 m1m2 m1m2 VCC VCC m1m2
+ VCC VCC VCC m1m2 bias1 m1m2 bias1 bias1 VCC bias1 VCC VCC bias1 VCC bias1 VCC m1m2
+ VCC m1m2 m1m2 bias1 bias1 VCC bias1 bias1 VCC bias1 VCC m1m2 m1m2 VCC bias1 bias1
+ VCC VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC VCC VCC bias1 m1m2 m1m2 bias1 m1m2 bias1
+ VCC VCC VCC VCC bias1 m1m2 m1m2 VCC bias1 bias1 VCC VCC bias1 VCC VCC m1m2 bias1
+ VCC VCC VCC bias1 m1m2 bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC bias1 VCC bias1
+ m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC VCC VCC VCC m1m2 bias1 bias1 VCC m1m2 VCC
+ VCC VCC bias1 bias1 VCC VCC VCC VCC m1m2 m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC
+ m1m2 bias1 VCC VCC VCC bias1 bias1 VCC VCC m1m2 m1m2 bias1 m1m2 VCC VCC bias1 m1m2
+ VCC bias1 m1m2 m1m2 VCC VCC m1m2 VCC VCC m1m2 VCC bias1 m1m2 m1m2 bias1 m1m2 VCC
+ bias1 VCC VCC bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC m1m2 VCC VCC VCC bias1 VCC
+ m1m2 VCC bias1 m1m2 VCC m1m2 m1m2 m1m2 VCC bias1 m1m2 VCC VCC VCC VCC bias1 VCC
+ bias1 m1m2 VCC m1m2 VCC m1m2 VCC VCC VCC bias1 VCC bias1 bias1 m1m2 bias1 VCC VCC
+ VCC VCC VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC bias1 VCC m1m2 m1m2 VCC
+ m1m2 VCC VCC VCC m1m2 sky130_fd_pr__pfet_01v8_F76D73
XXM100_dummy_4 IB VCC dummy_100 IB dummy_100 VCC dummy_100 dummy_100 sky130_fd_pr__pfet_01v8_P2UXFR
XXM100_dummy_5 IB dummy_100 VCC dummy_100 sky130_fd_pr__pfet_01v8_C2U9V5
XXM3_dummy_3 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
XXM1 m1m2 m1m2 bias1 VCC bias1 m1m2 VCC bias1 VCC VCC VCC bias1 m1m2 VCC VCC m1m2
+ VCC bias1 bias1 VCC VCC VCC bias1 m1m2 m1m2 m1m2 m1m2 bias1 VCC m1m2 VCC bias1 VCC
+ VCC VCC m1m2 m1m2 VCC bias1 VCC bias1 m1m2 bias1 VCC m1m2 VCC bias1 m1m2 VCC bias1
+ m1m2 VCC VCC VCC VCC VCC bias1 VCC VCC bias1 m1m2 m1m2 bias1 bias1 VCC VCC VCC m1m2
+ bias1 VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC VCC VCC VCC VCC m1m2 VCC m1m2 bias1
+ m1m2 bias1 VCC bias1 bias1 bias1 VCC VCC VCC bias1 m1m2 VCC m1m2 VCC bias1 m1m2
+ m1m2 VCC VCC bias1 VCC m1m2 m1m2 VCC bias1 VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC
+ m1m2 m1m2 VCC bias1 VCC VCC m1m2 VCC bias1 bias1 VCC VCC m1m2 VCC bias1 m1m2 VCC
+ m1m2 bias1 VCC VCC VCC m1m2 m1m2 VCC VCC VCC VCC VCC bias1 bias1 m1m2 m1m2 VCC m1m2
+ VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 bias1 VCC VCC m1m2 m1m2 m1m2 VCC VCC m1m2
+ VCC VCC VCC m1m2 bias1 m1m2 bias1 bias1 VCC bias1 VCC VCC bias1 VCC bias1 VCC m1m2
+ VCC m1m2 m1m2 bias1 bias1 VCC bias1 bias1 VCC bias1 VCC m1m2 m1m2 VCC bias1 bias1
+ VCC VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC VCC VCC bias1 m1m2 m1m2 bias1 m1m2 bias1
+ VCC VCC VCC VCC bias1 m1m2 m1m2 VCC bias1 bias1 VCC VCC bias1 VCC VCC m1m2 bias1
+ VCC VCC VCC bias1 m1m2 bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC bias1 VCC bias1
+ m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC VCC VCC VCC m1m2 bias1 bias1 VCC m1m2 VCC
+ VCC VCC bias1 bias1 VCC VCC VCC VCC m1m2 m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC
+ m1m2 bias1 VCC VCC VCC bias1 bias1 VCC VCC m1m2 m1m2 bias1 m1m2 VCC VCC bias1 m1m2
+ VCC bias1 m1m2 m1m2 VCC VCC m1m2 VCC VCC m1m2 VCC bias1 m1m2 m1m2 bias1 m1m2 VCC
+ bias1 VCC VCC bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC m1m2 VCC VCC VCC bias1 VCC
+ m1m2 VCC bias1 m1m2 VCC m1m2 m1m2 m1m2 VCC bias1 m1m2 VCC VCC VCC VCC bias1 VCC
+ bias1 m1m2 VCC m1m2 VCC m1m2 VCC VCC VCC bias1 VCC bias1 bias1 m1m2 bias1 VCC VCC
+ VCC VCC VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC bias1 VCC m1m2 m1m2 VCC
+ m1m2 VCC VCC VCC m1m2 sky130_fd_pr__pfet_01v8_F76D73
XXM100_dummy_6 IB dummy_100 VCC dummy_100 sky130_fd_pr__pfet_01v8_C2U9V5
XXM3_dummy_4 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
Xsky130_fd_pr__nfet_01v8_QP5WRD_0 bias1 bias1 VB_B bias1 VB_B VB_B VB_B VB_B m3m4
+ m3m4 m3m4 m3m4 bias1 bias1 VB_B bias1 bias1 VB_B bias1 bias1 m3m4 VB_B m3m4 m3m4
+ m3m4 m3m4 m3m4 VB_B VB_B bias1 bias1 VB_B bias1 VB_B bias1 VB_B VB_B m3m4 VB_B m3m4
+ m3m4 m3m4 m3m4 bias1 bias1 VSS sky130_fd_pr__nfet_01v8_QP5WRD
XXM2 bias1 VB_A m1m2 bias1 VB_A m1m2 VCC VCC m1m2 m1m2 m1m2 VB_A VCC m1m2 VCC bias1
+ VCC VCC VB_A bias1 VCC VB_A bias1 bias1 VB_A VB_A m1m2 VB_A m1m2 m1m2 bias1 m1m2
+ VCC m1m2 VCC VCC bias1 bias1 VCC bias1 bias1 bias1 VB_A VB_A VB_A VCC m1m2 VB_A
+ VCC VB_A m1m2 VCC VB_A m1m2 VCC VB_A m1m2 bias1 bias1 bias1 sky130_fd_pr__pfet_01v8_UDM5A5
XXM100_dummy_7 IB dummy_100 VCC dummy_100 sky130_fd_pr__pfet_01v8_C2U9V5
XXM4_dummy_10 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM8_1 VSS bias21 bias21 VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM3 m3m4 m3m4 VB_B m3m4 VB_B VB_B VB_B VB_B bias1 bias1 bias1 bias1 m3m4 m3m4 VB_B
+ m3m4 m3m4 VB_B m3m4 m3m4 bias1 VB_B bias1 bias1 bias1 bias1 bias1 VB_B VB_B m3m4
+ m3m4 VB_B m3m4 VB_B m3m4 VB_B VB_B bias1 VB_B bias1 bias1 bias1 bias1 m3m4 m3m4
+ VSS sky130_fd_pr__nfet_01v8_QP5WRD
XXM100_dummy_8 IB dummy_100 VCC dummy_100 sky130_fd_pr__pfet_01v8_C2U9V5
XXM3_dummy_6 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
XXM4 VSS m3m4 bias3 VSS sky130_fd_pr__nfet_01v8_3ZAA45
XXM100_dummy_9 IB dummy_100 VCC dummy_100 sky130_fd_pr__pfet_01v8_C2U9V5
XXM3_dummy_7 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
XXM8_3 VSS bias21 bias21 VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM5 VCC IN_M IN_M m1_44990_37960# VCC VCC bias3 bias3 bias3 m1_44990_37960# IN_M
+ m1_44990_37960# bias3 m1_44990_37960# IN_M bias3 m1_44990_37960# VCC IN_M IN_M m1_44990_37960#
+ VCC IN_M IN_M IN_M VCC VCC VCC IN_M IN_M IN_M bias3 bias3 bias3 m1_44990_37960#
+ IN_M VCC m1_44990_37960# bias3 m1_44990_37960# bias3 IN_M VCC m1_44990_37960# bias3
+ VCC m1_44990_37960# VCC VCC bias3 m1_44990_37960# bias3 m1_44990_37960# m1_44990_37960#
+ bias3 m1_44990_37960# VCC bias3 IN_M VCC sky130_fd_pr__pfet_01v8_7DHACV
XXM3_dummy_8 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
XXM6 bias3 bias3 VSS VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM6_1 bias3 bias3 VSS VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM3_dummy_9 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
Xsky130_fd_pr__pfet_01v8_SKU9VM_0 VB_A dummy_2 VCC dummy_2 sky130_fd_pr__pfet_01v8_SKU9VM
XXM7 VCC IN_P IN_P bias21 VCC VCC m1_44990_37960# m1_44990_37960# m1_44990_37960#
+ bias21 IN_P bias21 m1_44990_37960# bias21 IN_P m1_44990_37960# bias21 VCC IN_P IN_P
+ bias21 VCC IN_P IN_P IN_P VCC VCC VCC IN_P IN_P IN_P m1_44990_37960# m1_44990_37960#
+ m1_44990_37960# bias21 IN_P VCC bias21 m1_44990_37960# bias21 m1_44990_37960# IN_P
+ VCC bias21 m1_44990_37960# VCC bias21 VCC VCC m1_44990_37960# bias21 m1_44990_37960#
+ bias21 bias21 m1_44990_37960# bias21 VCC m1_44990_37960# IN_P VCC sky130_fd_pr__pfet_01v8_7DHACV
XXM6_2 bias3 bias3 VSS VSS sky130_fd_pr__nfet_01v8_VT3ZQW
Xsky130_fd_pr__pfet_01v8_E769TZ_0 dummy_9 dummy_9 bias1 VCC bias1 dummy_9 dummy_9
+ bias1 VCC VCC dummy_9 bias1 dummy_9 VCC VCC dummy_9 dummy_9 dummy_9 bias1 bias1
+ VCC VCC dummy_9 bias1 dummy_9 dummy_9 dummy_9 dummy_9 bias1 VCC dummy_9 dummy_9
+ bias1 VCC dummy_9 dummy_9 dummy_9 dummy_9 VCC bias1 VCC bias1 dummy_9 bias1 dummy_9
+ dummy_9 dummy_9 bias1 dummy_9 dummy_9 bias1 dummy_9 bias1 VCC VCC dummy_9 VCC VCC
+ bias1 dummy_9 dummy_9 bias1 dummy_9 dummy_9 bias1 bias1 VCC VCC dummy_9 dummy_9
+ bias1 dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1 dummy_9 VCC VCC dummy_9 VCC VCC
+ dummy_9 VCC dummy_9 bias1 dummy_9 bias1 dummy_9 bias1 bias1 bias1 VCC dummy_9 VCC
+ bias1 dummy_9 dummy_9 dummy_9 dummy_9 bias1 dummy_9 dummy_9 VCC bias1 VCC VCC dummy_9
+ dummy_9 dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1 VCC bias1 dummy_9 VCC dummy_9
+ dummy_9 dummy_9 VCC bias1 VCC dummy_9 dummy_9 dummy_9 bias1 bias1 dummy_9 dummy_9
+ dummy_9 dummy_9 VCC bias1 dummy_9 VCC dummy_9 bias1 VCC dummy_9 VCC dummy_9 dummy_9
+ dummy_9 VCC VCC dummy_9 VCC VCC bias1 bias1 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9
+ dummy_9 dummy_9 VCC VCC dummy_9 dummy_9 bias1 dummy_9 dummy_9 bias1 VCC dummy_9
+ dummy_9 dummy_9 dummy_9 VCC dummy_9 dummy_9 dummy_9 VCC VCC dummy_9 bias1 dummy_9
+ bias1 bias1 dummy_9 bias1 VCC dummy_9 bias1 VCC bias1 VCC dummy_9 VCC dummy_9 dummy_9
+ bias1 bias1 dummy_9 bias1 bias1 VCC bias1 dummy_9 dummy_9 dummy_9 VCC bias1 bias1
+ VCC VCC dummy_9 dummy_9 bias1 dummy_9 bias1 dummy_9 dummy_9 VCC bias1 dummy_9 bias1
+ dummy_9 dummy_9 bias1 dummy_9 bias1 VCC dummy_9 dummy_9 dummy_9 bias1 dummy_9 dummy_9
+ dummy_9 bias1 bias1 dummy_9 dummy_9 bias1 VCC dummy_9 dummy_9 bias1 VCC VCC dummy_9
+ bias1 dummy_9 bias1 dummy_9 bias1 VCC dummy_9 bias1 VCC dummy_9 dummy_9 bias1 dummy_9
+ bias1 dummy_9 dummy_9 VCC VCC VCC dummy_9 bias1 VCC VCC VCC dummy_9 dummy_9 dummy_9
+ bias1 bias1 dummy_9 dummy_9 VCC VCC VCC bias1 bias1 dummy_9 dummy_9 VCC VCC dummy_9
+ dummy_9 dummy_9 VCC VCC VCC VCC bias1 VCC VCC dummy_9 bias1 dummy_9 dummy_9 dummy_9
+ bias1 bias1 dummy_9 dummy_9 dummy_9 dummy_9 bias1 dummy_9 VCC VCC dummy_9 bias1
+ dummy_9 dummy_9 bias1 dummy_9 dummy_9 VCC VCC dummy_9 dummy_9 VCC dummy_9 dummy_9
+ bias1 dummy_9 dummy_9 bias1 dummy_9 dummy_9 bias1 dummy_9 VCC bias1 dummy_9 bias1
+ VCC dummy_9 bias1 VCC dummy_9 dummy_9 dummy_9 VCC VCC dummy_9 bias1 VCC dummy_9
+ dummy_9 bias1 dummy_9 VCC dummy_9 dummy_9 dummy_9 VCC bias1 dummy_9 dummy_9 VCC
+ VCC dummy_9 bias1 dummy_9 bias1 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9 VCC VCC
+ dummy_9 bias1 dummy_9 bias1 bias1 dummy_9 bias1 dummy_9 dummy_9 VCC VCC VCC dummy_9
+ dummy_9 dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1 VCC VCC bias1 dummy_9 dummy_9
+ dummy_9 VCC dummy_9 VCC VCC dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_E769TZ
XXM8 VSS bias21 bias21 VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM6_3 bias3 bias3 VSS VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM2_dummy_2 dummy_2 dummy_2 VB_A VB_A dummy_2 dummy_2 VB_A dummy_2 VCC VCC dummy_2
+ dummy_2 dummy_2 VB_A VCC dummy_2 dummy_2 VCC dummy_2 VCC VCC VB_A dummy_2 VCC VB_A
+ dummy_2 VCC dummy_2 VB_A VB_A dummy_2 VB_A dummy_2 dummy_2 dummy_2 dummy_2 dummy_2
+ VCC dummy_2 VCC VCC dummy_2 dummy_2 VCC dummy_2 dummy_2 dummy_2 VB_A VB_A VB_A VCC
+ dummy_2 VB_A VB_A VCC VB_A dummy_2 VCC VB_A dummy_2 VCC dummy_2 VB_A dummy_2 dummy_2
+ VCC dummy_2 dummy_2 sky130_fd_pr__pfet_01v8_UDMRD5
Xsky130_fd_pr__pfet_01v8_RRU5GE_0 IB VCC m1_44990_37960# VCC VCC IB VCC IB VCC VCC
+ m1_44990_37960# m1_44990_37960# sky130_fd_pr__pfet_01v8_RRU5GE
XXM9 VCC VCC bias1 VCC bias1 VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC m9m10 VCC
+ m9m10 bias1 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC m9m10 bias1
+ VCC m9m10 m9m10 VCC VCC VCC bias1 VCC bias1 VCC bias1 m9m10 VCC m9m10 bias1 VCC
+ m9m10 bias1 VCC VCC VCC m9m10 VCC VCC bias1 m9m10 m9m10 bias1 VCC VCC bias1 bias1
+ VCC VCC m9m10 VCC bias1 m9m10 bias1 m9m10 VCC m9m10 bias1 VCC VCC VCC m9m10 VCC
+ VCC VCC VCC VCC bias1 VCC bias1 m9m10 bias1 bias1 bias1 VCC m9m10 VCC bias1 VCC
+ m9m10 VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC VCC m9m10 bias1 m9m10 VCC VCC
+ bias1 VCC bias1 m9m10 VCC VCC VCC VCC bias1 VCC m9m10 VCC m9m10 bias1 bias1 m9m10
+ m9m10 VCC VCC bias1 VCC VCC VCC bias1 VCC m9m10 m9m10 VCC VCC VCC VCC m9m10 VCC
+ VCC bias1 bias1 VCC VCC m9m10 VCC m9m10 m9m10 VCC VCC VCC m9m10 bias1 m9m10 VCC
+ bias1 VCC m9m10 VCC VCC VCC VCC m9m10 VCC m9m10 VCC VCC VCC bias1 VCC bias1 bias1
+ m9m10 bias1 VCC m9m10 bias1 VCC bias1 VCC VCC VCC VCC VCC bias1 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC bias1 m9m10 bias1
+ m9m10 m9m10 VCC m9m10 bias1 VCC VCC bias1 VCC bias1 VCC m9m10 m9m10 m9m10 bias1
+ VCC VCC m9m10 bias1 bias1 m9m10 m9m10 bias1 VCC m9m10 VCC bias1 VCC VCC m9m10 bias1
+ VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 bias1 m9m10 bias1 VCC VCC
+ VCC VCC VCC m9m10 bias1 VCC VCC VCC m9m10 m9m10 VCC bias1 bias1 m9m10 VCC VCC VCC
+ VCC bias1 bias1 m9m10 m9m10 VCC VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC VCC
+ bias1 m9m10 m9m10 m9m10 bias1 bias1 m9m10 m9m10 VCC VCC bias1 VCC VCC VCC bias1
+ VCC m9m10 bias1 VCC VCC VCC VCC VCC m9m10 VCC VCC m9m10 bias1 VCC VCC bias1 VCC
+ m9m10 bias1 m9m10 VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 VCC VCC
+ VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC VCC VCC bias1 VCC m9m10 VCC
+ VCC m9m10 bias1 m9m10 bias1 VCC m9m10 VCC m9m10 VCC VCC VCC m9m10 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 m9m10 VCC VCC VCC m9m10 m9m10 m9m10 bias1 m9m10 m9m10 VCC
+ bias1 VCC VCC bias1 m9m10 VCC VCC VCC VCC VCC VCC m9m10 VCC sky130_fd_pr__pfet_01v8_F76D73
XXM2_dummy_3 VB_A dummy_2 VCC dummy_2 sky130_fd_pr__pfet_01v8_SKU9VM
Xsky130_fd_pr__pfet_01v8_C2U9V5_0 IB dummy_100 VCC dummy_100 sky130_fd_pr__pfet_01v8_C2U9V5
XXM2_dummy_4 VB_A dummy_2 VCC dummy_2 sky130_fd_pr__pfet_01v8_SKU9VM
Xsky130_fd_pr__nfet_01v8_AH5E2K_0 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
XXM2_dummy_5 VB_A dummy_2 VCC dummy_2 sky130_fd_pr__pfet_01v8_SKU9VM
XXM2_dummy_6 VB_A dummy_2 VCC dummy_2 sky130_fd_pr__pfet_01v8_SKU9VM
XXM2_1 m1m2 VB_A bias1 m1m2 VB_A bias1 VCC VCC bias1 bias1 bias1 VB_A VCC bias1 VCC
+ m1m2 VCC VCC VB_A m1m2 VCC VB_A m1m2 m1m2 VB_A VB_A bias1 VB_A bias1 bias1 m1m2
+ bias1 VCC bias1 VCC VCC m1m2 m1m2 VCC m1m2 m1m2 m1m2 VB_A VB_A VB_A VCC bias1 VB_A
+ VCC VB_A bias1 VCC VB_A bias1 VCC VB_A bias1 m1m2 m1m2 m1m2 sky130_fd_pr__pfet_01v8_UDM5A5
Xsky130_fd_pr__nfet_01v8_3ZAA45_0 m11m12 VSS bias21 VSS sky130_fd_pr__nfet_01v8_3ZAA45
XXM3_dummy_10 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
Xsky130_fd_pr__nfet_01v8_MHE452_0 dummy_4 bias3 dummy_4 dummy_4 bias3 dummy_4 bias3
+ dummy_4 bias3 dummy_4 dummy_4 dummy_4 dummy_4 dummy_4 bias3 dummy_4 dummy_4 bias3
+ VSS sky130_fd_pr__nfet_01v8_MHE452
XXM2_dummy_7 VB_A dummy_2 VCC dummy_2 sky130_fd_pr__pfet_01v8_SKU9VM
Xsky130_fd_pr__pfet_01v8_F76D73_0 m1m2 m1m2 bias1 VCC bias1 m1m2 VCC bias1 VCC VCC
+ VCC bias1 m1m2 VCC VCC m1m2 VCC bias1 bias1 VCC VCC VCC bias1 m1m2 m1m2 m1m2 m1m2
+ bias1 VCC m1m2 VCC bias1 VCC VCC VCC m1m2 m1m2 VCC bias1 VCC bias1 m1m2 bias1 VCC
+ m1m2 VCC bias1 m1m2 VCC bias1 m1m2 VCC VCC VCC VCC VCC bias1 VCC VCC bias1 m1m2
+ m1m2 bias1 bias1 VCC VCC VCC m1m2 bias1 VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC VCC
+ VCC VCC VCC m1m2 VCC m1m2 bias1 m1m2 bias1 VCC bias1 bias1 bias1 VCC VCC VCC bias1
+ m1m2 VCC m1m2 VCC bias1 m1m2 m1m2 VCC VCC bias1 VCC m1m2 m1m2 VCC bias1 VCC m1m2
+ m1m2 bias1 VCC bias1 VCC VCC m1m2 m1m2 VCC bias1 VCC VCC m1m2 VCC bias1 bias1 VCC
+ VCC m1m2 VCC bias1 m1m2 VCC m1m2 bias1 VCC VCC VCC m1m2 m1m2 VCC VCC VCC VCC VCC
+ bias1 bias1 m1m2 m1m2 VCC m1m2 VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 bias1 VCC
+ VCC m1m2 m1m2 m1m2 VCC VCC m1m2 VCC VCC VCC m1m2 bias1 m1m2 bias1 bias1 VCC bias1
+ VCC VCC bias1 VCC bias1 VCC m1m2 VCC m1m2 m1m2 bias1 bias1 VCC bias1 bias1 VCC bias1
+ VCC m1m2 m1m2 VCC bias1 bias1 VCC VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC VCC VCC
+ bias1 m1m2 m1m2 bias1 m1m2 bias1 VCC VCC VCC VCC bias1 m1m2 m1m2 VCC bias1 bias1
+ VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC VCC bias1 m1m2 bias1 VCC bias1 VCC VCC
+ bias1 VCC VCC VCC bias1 VCC bias1 m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC VCC VCC
+ VCC m1m2 bias1 bias1 VCC m1m2 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC m1m2 m1m2
+ m1m2 VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC VCC bias1 bias1 VCC VCC m1m2
+ m1m2 bias1 m1m2 VCC VCC bias1 m1m2 VCC bias1 m1m2 m1m2 VCC VCC m1m2 VCC VCC m1m2
+ VCC bias1 m1m2 m1m2 bias1 m1m2 VCC bias1 VCC VCC bias1 VCC bias1 VCC VCC bias1 VCC
+ VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC m1m2 m1m2 m1m2 VCC bias1
+ m1m2 VCC VCC VCC VCC bias1 VCC bias1 m1m2 VCC m1m2 VCC m1m2 VCC VCC VCC bias1 VCC
+ bias1 bias1 m1m2 bias1 VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1
+ VCC VCC bias1 VCC m1m2 m1m2 VCC m1m2 VCC VCC VCC m1m2 sky130_fd_pr__pfet_01v8_F76D73
Xsky130_fd_pr__pfet_01v8_UDM5A5_0 m9m10 VB_A OUT m9m10 VB_A OUT VCC VCC OUT OUT OUT
+ VB_A VCC OUT VCC m9m10 VCC VCC VB_A m9m10 VCC VB_A m9m10 m9m10 VB_A VB_A OUT VB_A
+ OUT OUT m9m10 OUT VCC OUT VCC VCC m9m10 m9m10 VCC m9m10 m9m10 m9m10 VB_A VB_A VB_A
+ VCC OUT VB_A VCC VB_A OUT VCC VB_A OUT VCC VB_A OUT m9m10 m9m10 m9m10 sky130_fd_pr__pfet_01v8_UDM5A5
XXM9_dummy_1 dummy_9 dummy_9 bias1 VCC bias1 dummy_9 dummy_9 bias1 VCC VCC dummy_9
+ bias1 dummy_9 VCC VCC dummy_9 dummy_9 dummy_9 bias1 bias1 VCC VCC dummy_9 bias1
+ dummy_9 dummy_9 dummy_9 dummy_9 bias1 VCC dummy_9 dummy_9 bias1 VCC dummy_9 dummy_9
+ dummy_9 dummy_9 VCC bias1 VCC bias1 dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1
+ dummy_9 dummy_9 bias1 dummy_9 bias1 VCC VCC dummy_9 VCC VCC bias1 dummy_9 dummy_9
+ bias1 dummy_9 dummy_9 bias1 bias1 VCC VCC dummy_9 dummy_9 bias1 dummy_9 bias1 dummy_9
+ dummy_9 dummy_9 bias1 dummy_9 VCC VCC dummy_9 VCC VCC dummy_9 VCC dummy_9 bias1
+ dummy_9 bias1 dummy_9 bias1 bias1 bias1 VCC dummy_9 VCC bias1 dummy_9 dummy_9 dummy_9
+ dummy_9 bias1 dummy_9 dummy_9 VCC bias1 VCC VCC dummy_9 dummy_9 dummy_9 bias1 dummy_9
+ dummy_9 dummy_9 bias1 VCC bias1 dummy_9 VCC dummy_9 dummy_9 dummy_9 VCC bias1 VCC
+ dummy_9 dummy_9 dummy_9 bias1 bias1 dummy_9 dummy_9 dummy_9 dummy_9 VCC bias1 dummy_9
+ VCC dummy_9 bias1 VCC dummy_9 VCC dummy_9 dummy_9 dummy_9 VCC VCC dummy_9 VCC VCC
+ bias1 bias1 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9 VCC VCC dummy_9
+ dummy_9 bias1 dummy_9 dummy_9 bias1 VCC dummy_9 dummy_9 dummy_9 dummy_9 VCC dummy_9
+ dummy_9 dummy_9 VCC VCC dummy_9 bias1 dummy_9 bias1 bias1 dummy_9 bias1 VCC dummy_9
+ bias1 VCC bias1 VCC dummy_9 VCC dummy_9 dummy_9 bias1 bias1 dummy_9 bias1 bias1
+ VCC bias1 dummy_9 dummy_9 dummy_9 VCC bias1 bias1 VCC VCC dummy_9 dummy_9 bias1
+ dummy_9 bias1 dummy_9 dummy_9 VCC bias1 dummy_9 bias1 dummy_9 dummy_9 bias1 dummy_9
+ bias1 VCC dummy_9 dummy_9 dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1 bias1 dummy_9
+ dummy_9 bias1 VCC dummy_9 dummy_9 bias1 VCC VCC dummy_9 bias1 dummy_9 bias1 dummy_9
+ bias1 VCC dummy_9 bias1 VCC dummy_9 dummy_9 bias1 dummy_9 bias1 dummy_9 dummy_9
+ VCC VCC VCC dummy_9 bias1 VCC VCC VCC dummy_9 dummy_9 dummy_9 bias1 bias1 dummy_9
+ dummy_9 VCC VCC VCC bias1 bias1 dummy_9 dummy_9 VCC VCC dummy_9 dummy_9 dummy_9
+ VCC VCC VCC VCC bias1 VCC VCC dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1 bias1
+ dummy_9 dummy_9 dummy_9 dummy_9 bias1 dummy_9 VCC VCC dummy_9 bias1 dummy_9 dummy_9
+ bias1 dummy_9 dummy_9 VCC VCC dummy_9 dummy_9 VCC dummy_9 dummy_9 bias1 dummy_9
+ dummy_9 bias1 dummy_9 dummy_9 bias1 dummy_9 VCC bias1 dummy_9 bias1 VCC dummy_9
+ bias1 VCC dummy_9 dummy_9 dummy_9 VCC VCC dummy_9 bias1 VCC dummy_9 dummy_9 bias1
+ dummy_9 VCC dummy_9 dummy_9 dummy_9 VCC bias1 dummy_9 dummy_9 VCC VCC dummy_9 bias1
+ dummy_9 bias1 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9 VCC VCC dummy_9 bias1 dummy_9
+ bias1 bias1 dummy_9 bias1 dummy_9 dummy_9 VCC VCC VCC dummy_9 dummy_9 dummy_9 bias1
+ dummy_9 dummy_9 dummy_9 bias1 VCC VCC bias1 dummy_9 dummy_9 dummy_9 VCC dummy_9
+ VCC VCC dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_E769TZ
XXM2_dummy_9 VB_A dummy_2 VCC dummy_2 sky130_fd_pr__pfet_01v8_SKU9VM
XXM9_dummy_3 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_SLZ774
XXM9_dummy_4 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_dummy_5 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
Xsky130_fd_pr__pfet_01v8_UDMRD5_0 dummy_2 dummy_2 VB_A VB_A dummy_2 dummy_2 VB_A dummy_2
+ VCC VCC dummy_2 dummy_2 dummy_2 VB_A VCC dummy_2 dummy_2 VCC dummy_2 VCC VCC VB_A
+ dummy_2 VCC VB_A dummy_2 VCC dummy_2 VB_A VB_A dummy_2 VB_A dummy_2 dummy_2 dummy_2
+ dummy_2 dummy_2 VCC dummy_2 VCC VCC dummy_2 dummy_2 VCC dummy_2 dummy_2 dummy_2
+ VB_A VB_A VB_A VCC dummy_2 VB_A VB_A VCC VB_A dummy_2 VCC VB_A dummy_2 VCC dummy_2
+ VB_A dummy_2 dummy_2 VCC dummy_2 dummy_2 sky130_fd_pr__pfet_01v8_UDMRD5
XXM9_dummy_20 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_1 VCC VCC bias1 VCC bias1 VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC m9m10 VCC
+ m9m10 bias1 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC m9m10 bias1
+ VCC m9m10 m9m10 VCC VCC VCC bias1 VCC bias1 VCC bias1 m9m10 VCC m9m10 bias1 VCC
+ m9m10 bias1 VCC VCC VCC m9m10 VCC VCC bias1 m9m10 m9m10 bias1 VCC VCC bias1 bias1
+ VCC VCC m9m10 VCC bias1 m9m10 bias1 m9m10 VCC m9m10 bias1 VCC VCC VCC m9m10 VCC
+ VCC VCC VCC VCC bias1 VCC bias1 m9m10 bias1 bias1 bias1 VCC m9m10 VCC bias1 VCC
+ m9m10 VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC VCC m9m10 bias1 m9m10 VCC VCC
+ bias1 VCC bias1 m9m10 VCC VCC VCC VCC bias1 VCC m9m10 VCC m9m10 bias1 bias1 m9m10
+ m9m10 VCC VCC bias1 VCC VCC VCC bias1 VCC m9m10 m9m10 VCC VCC VCC VCC m9m10 VCC
+ VCC bias1 bias1 VCC VCC m9m10 VCC m9m10 m9m10 VCC VCC VCC m9m10 bias1 m9m10 VCC
+ bias1 VCC m9m10 VCC VCC VCC VCC m9m10 VCC m9m10 VCC VCC VCC bias1 VCC bias1 bias1
+ m9m10 bias1 VCC m9m10 bias1 VCC bias1 VCC VCC VCC VCC VCC bias1 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC bias1 m9m10 bias1
+ m9m10 m9m10 VCC m9m10 bias1 VCC VCC bias1 VCC bias1 VCC m9m10 m9m10 m9m10 bias1
+ VCC VCC m9m10 bias1 bias1 m9m10 m9m10 bias1 VCC m9m10 VCC bias1 VCC VCC m9m10 bias1
+ VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 bias1 m9m10 bias1 VCC VCC
+ VCC VCC VCC m9m10 bias1 VCC VCC VCC m9m10 m9m10 VCC bias1 bias1 m9m10 VCC VCC VCC
+ VCC bias1 bias1 m9m10 m9m10 VCC VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC VCC
+ bias1 m9m10 m9m10 m9m10 bias1 bias1 m9m10 m9m10 VCC VCC bias1 VCC VCC VCC bias1
+ VCC m9m10 bias1 VCC VCC VCC VCC VCC m9m10 VCC VCC m9m10 bias1 VCC VCC bias1 VCC
+ m9m10 bias1 m9m10 VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 VCC VCC
+ VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC VCC VCC bias1 VCC m9m10 VCC
+ VCC m9m10 bias1 m9m10 bias1 VCC m9m10 VCC m9m10 VCC VCC VCC m9m10 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 m9m10 VCC VCC VCC m9m10 m9m10 m9m10 bias1 m9m10 m9m10 VCC
+ bias1 VCC VCC bias1 m9m10 VCC VCC VCC VCC VCC VCC m9m10 VCC sky130_fd_pr__pfet_01v8_F76D73
XXM9_dummy_6 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_dummy_10 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_2 VCC VCC bias1 VCC bias1 VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC m9m10 VCC
+ m9m10 bias1 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC m9m10 bias1
+ VCC m9m10 m9m10 VCC VCC VCC bias1 VCC bias1 VCC bias1 m9m10 VCC m9m10 bias1 VCC
+ m9m10 bias1 VCC VCC VCC m9m10 VCC VCC bias1 m9m10 m9m10 bias1 VCC VCC bias1 bias1
+ VCC VCC m9m10 VCC bias1 m9m10 bias1 m9m10 VCC m9m10 bias1 VCC VCC VCC m9m10 VCC
+ VCC VCC VCC VCC bias1 VCC bias1 m9m10 bias1 bias1 bias1 VCC m9m10 VCC bias1 VCC
+ m9m10 VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC VCC m9m10 bias1 m9m10 VCC VCC
+ bias1 VCC bias1 m9m10 VCC VCC VCC VCC bias1 VCC m9m10 VCC m9m10 bias1 bias1 m9m10
+ m9m10 VCC VCC bias1 VCC VCC VCC bias1 VCC m9m10 m9m10 VCC VCC VCC VCC m9m10 VCC
+ VCC bias1 bias1 VCC VCC m9m10 VCC m9m10 m9m10 VCC VCC VCC m9m10 bias1 m9m10 VCC
+ bias1 VCC m9m10 VCC VCC VCC VCC m9m10 VCC m9m10 VCC VCC VCC bias1 VCC bias1 bias1
+ m9m10 bias1 VCC m9m10 bias1 VCC bias1 VCC VCC VCC VCC VCC bias1 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC bias1 m9m10 bias1
+ m9m10 m9m10 VCC m9m10 bias1 VCC VCC bias1 VCC bias1 VCC m9m10 m9m10 m9m10 bias1
+ VCC VCC m9m10 bias1 bias1 m9m10 m9m10 bias1 VCC m9m10 VCC bias1 VCC VCC m9m10 bias1
+ VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 bias1 m9m10 bias1 VCC VCC
+ VCC VCC VCC m9m10 bias1 VCC VCC VCC m9m10 m9m10 VCC bias1 bias1 m9m10 VCC VCC VCC
+ VCC bias1 bias1 m9m10 m9m10 VCC VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC VCC
+ bias1 m9m10 m9m10 m9m10 bias1 bias1 m9m10 m9m10 VCC VCC bias1 VCC VCC VCC bias1
+ VCC m9m10 bias1 VCC VCC VCC VCC VCC m9m10 VCC VCC m9m10 bias1 VCC VCC bias1 VCC
+ m9m10 bias1 m9m10 VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 VCC VCC
+ VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC VCC VCC bias1 VCC m9m10 VCC
+ VCC m9m10 bias1 m9m10 bias1 VCC m9m10 VCC m9m10 VCC VCC VCC m9m10 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 m9m10 VCC VCC VCC m9m10 m9m10 m9m10 bias1 m9m10 m9m10 VCC
+ bias1 VCC VCC bias1 m9m10 VCC VCC VCC VCC VCC VCC m9m10 VCC sky130_fd_pr__pfet_01v8_F76D73
XXM9_dummy_7 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_dummy_22 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_dummy_11 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_3 VCC VCC bias1 VCC bias1 VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC m9m10 VCC
+ m9m10 bias1 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC m9m10 bias1
+ VCC m9m10 m9m10 VCC VCC VCC bias1 VCC bias1 VCC bias1 m9m10 VCC m9m10 bias1 VCC
+ m9m10 bias1 VCC VCC VCC m9m10 VCC VCC bias1 m9m10 m9m10 bias1 VCC VCC bias1 bias1
+ VCC VCC m9m10 VCC bias1 m9m10 bias1 m9m10 VCC m9m10 bias1 VCC VCC VCC m9m10 VCC
+ VCC VCC VCC VCC bias1 VCC bias1 m9m10 bias1 bias1 bias1 VCC m9m10 VCC bias1 VCC
+ m9m10 VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC VCC m9m10 bias1 m9m10 VCC VCC
+ bias1 VCC bias1 m9m10 VCC VCC VCC VCC bias1 VCC m9m10 VCC m9m10 bias1 bias1 m9m10
+ m9m10 VCC VCC bias1 VCC VCC VCC bias1 VCC m9m10 m9m10 VCC VCC VCC VCC m9m10 VCC
+ VCC bias1 bias1 VCC VCC m9m10 VCC m9m10 m9m10 VCC VCC VCC m9m10 bias1 m9m10 VCC
+ bias1 VCC m9m10 VCC VCC VCC VCC m9m10 VCC m9m10 VCC VCC VCC bias1 VCC bias1 bias1
+ m9m10 bias1 VCC m9m10 bias1 VCC bias1 VCC VCC VCC VCC VCC bias1 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC bias1 m9m10 bias1
+ m9m10 m9m10 VCC m9m10 bias1 VCC VCC bias1 VCC bias1 VCC m9m10 m9m10 m9m10 bias1
+ VCC VCC m9m10 bias1 bias1 m9m10 m9m10 bias1 VCC m9m10 VCC bias1 VCC VCC m9m10 bias1
+ VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 bias1 m9m10 bias1 VCC VCC
+ VCC VCC VCC m9m10 bias1 VCC VCC VCC m9m10 m9m10 VCC bias1 bias1 m9m10 VCC VCC VCC
+ VCC bias1 bias1 m9m10 m9m10 VCC VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC VCC
+ bias1 m9m10 m9m10 m9m10 bias1 bias1 m9m10 m9m10 VCC VCC bias1 VCC VCC VCC bias1
+ VCC m9m10 bias1 VCC VCC VCC VCC VCC m9m10 VCC VCC m9m10 bias1 VCC VCC bias1 VCC
+ m9m10 bias1 m9m10 VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 VCC VCC
+ VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC VCC VCC bias1 VCC m9m10 VCC
+ VCC m9m10 bias1 m9m10 bias1 VCC m9m10 VCC m9m10 VCC VCC VCC m9m10 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 m9m10 VCC VCC VCC m9m10 m9m10 m9m10 bias1 m9m10 m9m10 VCC
+ bias1 VCC VCC bias1 m9m10 VCC VCC VCC VCC VCC VCC m9m10 VCC sky130_fd_pr__pfet_01v8_F76D73
XXM11_1 OUT OUT VB_B OUT VB_B VB_B VB_B VB_B m11m12 m11m12 m11m12 m11m12 OUT OUT VB_B
+ OUT OUT VB_B OUT OUT m11m12 VB_B m11m12 m11m12 m11m12 m11m12 m11m12 VB_B VB_B OUT
+ OUT VB_B OUT VB_B OUT VB_B VB_B m11m12 VB_B m11m12 m11m12 m11m12 m11m12 OUT OUT
+ VSS sky130_fd_pr__nfet_01v8_QP5WRD
XXM9_dummy_8 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
Xsky130_fd_pr__nfet_01v8_SCE452_0 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM9_4 VCC VCC bias1 VCC bias1 VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC m9m10 VCC
+ m9m10 bias1 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC m9m10 bias1
+ VCC m9m10 m9m10 VCC VCC VCC bias1 VCC bias1 VCC bias1 m9m10 VCC m9m10 bias1 VCC
+ m9m10 bias1 VCC VCC VCC m9m10 VCC VCC bias1 m9m10 m9m10 bias1 VCC VCC bias1 bias1
+ VCC VCC m9m10 VCC bias1 m9m10 bias1 m9m10 VCC m9m10 bias1 VCC VCC VCC m9m10 VCC
+ VCC VCC VCC VCC bias1 VCC bias1 m9m10 bias1 bias1 bias1 VCC m9m10 VCC bias1 VCC
+ m9m10 VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC VCC m9m10 bias1 m9m10 VCC VCC
+ bias1 VCC bias1 m9m10 VCC VCC VCC VCC bias1 VCC m9m10 VCC m9m10 bias1 bias1 m9m10
+ m9m10 VCC VCC bias1 VCC VCC VCC bias1 VCC m9m10 m9m10 VCC VCC VCC VCC m9m10 VCC
+ VCC bias1 bias1 VCC VCC m9m10 VCC m9m10 m9m10 VCC VCC VCC m9m10 bias1 m9m10 VCC
+ bias1 VCC m9m10 VCC VCC VCC VCC m9m10 VCC m9m10 VCC VCC VCC bias1 VCC bias1 bias1
+ m9m10 bias1 VCC m9m10 bias1 VCC bias1 VCC VCC VCC VCC VCC bias1 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC bias1 m9m10 bias1
+ m9m10 m9m10 VCC m9m10 bias1 VCC VCC bias1 VCC bias1 VCC m9m10 m9m10 m9m10 bias1
+ VCC VCC m9m10 bias1 bias1 m9m10 m9m10 bias1 VCC m9m10 VCC bias1 VCC VCC m9m10 bias1
+ VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 bias1 m9m10 bias1 VCC VCC
+ VCC VCC VCC m9m10 bias1 VCC VCC VCC m9m10 m9m10 VCC bias1 bias1 m9m10 VCC VCC VCC
+ VCC bias1 bias1 m9m10 m9m10 VCC VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC VCC
+ bias1 m9m10 m9m10 m9m10 bias1 bias1 m9m10 m9m10 VCC VCC bias1 VCC VCC VCC bias1
+ VCC m9m10 bias1 VCC VCC VCC VCC VCC m9m10 VCC VCC m9m10 bias1 VCC VCC bias1 VCC
+ m9m10 bias1 m9m10 VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 VCC VCC
+ VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC VCC VCC bias1 VCC m9m10 VCC
+ VCC m9m10 bias1 m9m10 bias1 VCC m9m10 VCC m9m10 VCC VCC VCC m9m10 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 m9m10 VCC VCC VCC m9m10 m9m10 m9m10 bias1 m9m10 m9m10 VCC
+ bias1 VCC VCC bias1 m9m10 VCC VCC VCC VCC VCC VCC m9m10 VCC sky130_fd_pr__pfet_01v8_F76D73
XXM9_dummy_12 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM10 OUT VB_A m9m10 OUT VB_A m9m10 VCC VCC m9m10 m9m10 m9m10 VB_A VCC m9m10 VCC OUT
+ VCC VCC VB_A OUT VCC VB_A OUT OUT VB_A VB_A m9m10 VB_A m9m10 m9m10 OUT m9m10 VCC
+ m9m10 VCC VCC OUT OUT VCC OUT OUT OUT VB_A VB_A VB_A VCC m9m10 VB_A VCC VB_A m9m10
+ VCC VB_A m9m10 VCC VB_A m9m10 OUT OUT OUT sky130_fd_pr__pfet_01v8_UDM5A5
XXM9_dummy_9 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
Xsky130_fd_pr__pfet_01v8_7DHACV_0 VCC IN_P IN_P m1_44990_37960# VCC VCC bias21 bias21
+ bias21 m1_44990_37960# IN_P m1_44990_37960# bias21 m1_44990_37960# IN_P bias21 m1_44990_37960#
+ VCC IN_P IN_P m1_44990_37960# VCC IN_P IN_P IN_P VCC VCC VCC IN_P IN_P IN_P bias21
+ bias21 bias21 m1_44990_37960# IN_P VCC m1_44990_37960# bias21 m1_44990_37960# bias21
+ IN_P VCC m1_44990_37960# bias21 VCC m1_44990_37960# VCC VCC bias21 m1_44990_37960#
+ bias21 m1_44990_37960# m1_44990_37960# bias21 m1_44990_37960# VCC bias21 IN_P VCC
+ sky130_fd_pr__pfet_01v8_7DHACV
Xsky130_fd_pr__nfet_01v8_SCE452_1 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM9_dummy_13 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM100_1 IB VCC VCC m1_44990_37960# VCC IB m1_44990_37960# IB VCC m1_44990_37960#
+ VCC VCC sky130_fd_pr__pfet_01v8_RRU5GE
XXM11 m11m12 m11m12 VB_B m11m12 VB_B VB_B VB_B VB_B OUT OUT OUT OUT m11m12 m11m12
+ VB_B m11m12 m11m12 VB_B m11m12 m11m12 OUT VB_B OUT OUT OUT OUT OUT VB_B VB_B m11m12
+ m11m12 VB_B m11m12 VB_B m11m12 VB_B VB_B OUT VB_B OUT OUT OUT OUT m11m12 m11m12
+ VSS sky130_fd_pr__nfet_01v8_QP5WRD
XXM2_dummy_10 VB_A dummy_2 VCC dummy_2 sky130_fd_pr__pfet_01v8_SKU9VM
Xsky130_fd_pr__nfet_01v8_WK8VRD_0 VB_B dummy_3 dummy_3 dummy_3 VB_B dummy_3 VB_B VB_B
+ VB_B VB_B dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 VB_B dummy_3 dummy_3 dummy_3
+ VB_B dummy_3 dummy_3 dummy_3 VB_B dummy_3 dummy_3 dummy_3 dummy_3 VB_B dummy_3 dummy_3
+ VB_B VB_B dummy_3 dummy_3 VB_B dummy_3 VB_B dummy_3 VB_B VB_B dummy_3 VB_B dummy_3
+ dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 VSS sky130_fd_pr__nfet_01v8_WK8VRD
Xsky130_fd_pr__nfet_01v8_SCE452_2 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM9_dummy_14 VCC bias1 dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_ZLZ7XS
.ends

