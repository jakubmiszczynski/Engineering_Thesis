** sch_path: /home/kuba/project/SKY130_OpAmp/06_ParasiticsSim/opamp_cascode_dc_max_gain_mc.sch
**.subckt opamp_cascode_dc_max_gain_mc
Vcm net1 GND 0.985
.save i(vcm)
C1 out GND 1p m=1
Vdiff Vdiff GND 0
.save i(vdiff)
Ib IBIAS GND 45u
B1 Vp net1 v=v(Vdiff)
B2 net1 Vn v=v(Vdiff)
x1 Vp Vn VCC GND out VB_A VB_B IBIAS opamp_cascode
**** begin user architecture code


Vsupply VCC GND 1.8
VbiasA VB_A GND 0.2
VbiasB VB_B GND 1.1
.include ../opamp_cascode.spice
.control
  set wr_vecnames
  set wr_singlescale
  let mc_runs=5
  let run=1
  set curplot=new
  set final=$curplot
  setplot $final
  dowhile run <= mc_runs
    save all
    dc Vdiff -0.01 0.01 0.000001
    let dVout = deriv(v(out))
    meas dc maxGain max dVout
    set dt = $curplot
    setplot $final
    let dVout{$&run}={$dt}.v(dVout)
    let maxGain{$&run}={$dt}.maxGain
    setplot $dt
    reset
    let run = run + 1
  end
  setplot $final
  plot allv vs dc1.v(Vdiff) retraceplot
  set hcopydevtype = svg
  hardcopy dc_max_gain_mc.svg allv vs dc1.v(Vdiff)
.endc



.param mc_mm_switch=1
.param mc_pr_switch=0
.include ~/.volare/sky130A/libs.tech/ngspice/corners/tt.spice
.include ~/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include ~/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include ~/.volare/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
