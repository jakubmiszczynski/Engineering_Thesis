* NGSPICE file created from opamp_cascode.ext - technology: sky130A

.subckt opamp_cascode IN_P IN_M VCC VSS OUT VB_A VB_B IB
X0 m9m10.t499 bias1.t7 VCC.t1036 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1 VCC.t1035 bias1.t8 m1m2.t499 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X2 m3m4.t29 VB_B.t0 bias1.t2 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X3 dummy_9.t447 bias1.t9 dummy_9.t446 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X4 VCC.t1034 bias1.t10 m1m2.t498 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X5 dummy_9.t445 bias1.t11 dummy_9.t444 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X6 VCC.t1033 bias1.t12 m1m2.t497 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X7 m9m10.t498 bias1.t13 VCC.t1032 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X8 dummy_9.t443 bias1.t14 dummy_9.t442 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X9 m9m10.t497 bias1.t15 VCC.t1031 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X10 dummy_4.t39 bias3.t38 dummy_4.t38 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X11 VCC.t1030 bias1.t16 m1m2.t496 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X12 m9m10.t496 bias1.t17 VCC.t1029 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X13 dummy_9.t441 bias1.t18 dummy_9.t440 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X14 dummy_9.t439 bias1.t19 dummy_9.t438 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X15 m9m10.t495 bias1.t20 VCC.t1028 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X16 dummy_4.t37 bias3.t39 dummy_4.t36 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X17 m9m10.t494 bias1.t21 VCC.t1027 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X18 dummy_9.t437 bias1.t22 dummy_9.t436 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X19 VCC.t1026 bias1.t23 m1m2.t495 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X20 m9m10.t493 bias1.t24 VCC.t1025 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X21 m9m10.t492 bias1.t25 VCC.t1024 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X22 m1m2.t521 VB_A.t0 bias1.t6 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X23 dummy_9.t435 bias1.t26 dummy_9.t434 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X24 m9m10.t491 bias1.t27 VCC.t1023 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X25 m9m10.t490 bias1.t28 VCC.t1022 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X26 dummy_100.t39 IB.t8 dummy_100.t38 VCC.t7 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X27 VCC.t1021 bias1.t29 m1m2.t494 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X28 dummy_3.t83 VB_B.t1 dummy_3.t82 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X29 VCC.t1020 bias1.t30 m1m2.t493 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X30 m9m10.t489 bias1.t31 VCC.t1019 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X31 m9m10.t488 bias1.t32 VCC.t1018 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X32 dummy_9.t433 bias1.t33 dummy_9.t432 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X33 dummy_2.t83 VB_A.t1 dummy_2.t82 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X34 dummy_3.t81 VB_B.t2 dummy_3.t80 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X35 VCC.t1017 bias1.t34 m1m2.t492 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X36 m9m10.t487 bias1.t35 VCC.t1016 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X37 m9m10.t486 bias1.t36 VCC.t1015 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X38 m9m10.t485 bias1.t37 VCC.t1014 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X39 m9m10.t484 bias1.t38 VCC.t1013 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X40 VCC.t1012 bias1.t39 m1m2.t491 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X41 dummy_9.t431 bias1.t40 dummy_9.t430 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X42 VCC.t1011 bias1.t41 m1m2.t490 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X43 VCC.t1010 bias1.t42 m1m2.t489 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X44 m9m10.t483 bias1.t43 VCC.t976 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X45 dummy_100.t37 IB.t9 dummy_100.t36 VCC.t8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X46 m9m10.t482 bias1.t44 VCC.t1009 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X47 OUT.t29 VB_A.t2 m9m10.t522 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X48 m1m2.t519 VB_A.t3 bias1.t6 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X49 VCC.t1008 bias1.t45 m1m2.t488 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X50 m9m10.t481 bias1.t46 VCC.t986 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X51 VCC.t1007 bias1.t47 m1m2.t487 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X52 m9m10.t480 bias1.t48 VCC.t1006 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X53 dummy_9.t429 bias1.t49 dummy_9.t428 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X54 dummy_9.t427 bias1.t50 dummy_9.t426 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X55 VCC.t979 bias1.t51 m1m2.t486 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X56 dummy_4.t35 bias3.t40 dummy_4.t34 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X57 m9m10.t479 bias1.t52 VCC.t1005 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X58 dummy_2.t81 VB_A.t4 dummy_2.t80 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X59 VCC.t1004 bias1.t53 m1m2.t485 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X60 VCC.t978 bias1.t54 m1m2.t484 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X61 m9m10.t478 bias1.t55 VCC.t1003 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X62 m9m10.t477 bias1.t56 VCC.t985 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X63 dummy_9.t425 bias1.t57 dummy_9.t424 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X64 VCC.t977 bias1.t58 m1m2.t483 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X65 VCC.t981 bias1.t59 m1m2.t482 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X66 a_46836_49340.t45 IN_M.t0 bias3.t28 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X67 m9m10.t476 bias1.t60 VCC.t984 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X68 m9m10.t475 bias1.t61 VCC.t1002 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X69 VCC.t1001 bias1.t62 m1m2.t481 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X70 dummy_9.t423 bias1.t63 dummy_9.t422 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X71 m9m10.t474 bias1.t64 VCC.t1000 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X72 VCC.t980 bias1.t65 m1m2.t480 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X73 m9m10.t473 bias1.t66 VCC.t999 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X74 dummy_9.t421 bias1.t67 dummy_9.t420 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X75 m9m10.t472 bias1.t68 VCC.t998 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X76 dummy_9.t419 bias1.t69 dummy_9.t418 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X77 dummy_9.t417 bias1.t70 dummy_9.t416 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X78 m9m10.t471 bias1.t71 VCC.t997 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X79 VCC.t996 bias1.t72 m1m2.t479 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X80 m9m10.t470 bias1.t73 VCC.t995 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X81 m9m10.t469 bias1.t74 VCC.t994 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X82 VCC.t993 bias1.t75 m1m2.t478 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X83 m9m10.t468 bias1.t76 VCC.t992 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X84 VCC.t988 bias1.t77 m1m2.t477 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X85 m9m10.t467 bias1.t78 VCC.t991 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X86 dummy_9.t415 bias1.t57 dummy_9.t414 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X87 VCC.t990 bias1.t79 m1m2.t476 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X88 dummy_9.t413 bias1.t80 dummy_9.t412 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X89 m9m10.t466 bias1.t81 VCC.t989 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X90 VCC.t987 bias1.t82 m1m2.t475 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X91 dummy_9.t411 bias1.t83 dummy_9.t410 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X92 m3m4.t28 VB_B.t3 bias1.t2 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X93 dummy_9.t409 bias1.t84 dummy_9.t408 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X94 m9m10.t465 bias1.t85 VCC.t983 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X95 VCC.t982 bias1.t86 m1m2.t474 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X96 VCC.t975 bias1.t87 m1m2.t473 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X97 m9m10.t464 bias1.t88 VCC.t974 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X98 VCC.t973 bias1.t89 m1m2.t472 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X99 VCC.t972 bias1.t90 m1m2.t471 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X100 VCC.t971 bias1.t91 m1m2.t470 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X101 dummy_9.t407 bias1.t92 dummy_9.t406 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X102 VCC.t970 bias1.t93 m1m2.t469 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X103 bias21.t37 IN_P.t0 a_46836_49340.t54 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X104 m9m10.t521 VB_A.t5 OUT.t28 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X105 VCC.t969 bias1.t94 m1m2.t468 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X106 VCC.t968 bias1.t95 m1m2.t467 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X107 dummy_100.t35 IB.t10 dummy_100.t34 VCC.t8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X108 bias1.t6 VB_A.t6 m1m2.t515 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X109 m9m10.t463 bias1.t96 VCC.t967 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X110 VCC.t966 bias1.t97 m1m2.t466 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X111 VCC.t965 bias1.t98 m1m2.t465 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X112 m9m10.t462 bias1.t99 VCC.t964 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X113 dummy_9.t405 bias1.t100 dummy_9.t404 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X114 m9m10.t461 bias1.t101 VCC.t963 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X115 dummy_9.t403 bias1.t102 dummy_9.t402 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X116 m9m10.t460 bias1.t103 VCC.t962 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X117 VCC.t961 bias1.t104 m1m2.t464 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X118 m9m10.t459 bias1.t105 VCC.t960 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X119 dummy_9.t401 bias1.t106 dummy_9.t400 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X120 VCC.t959 bias1.t107 m1m2.t463 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X121 a_46836_49340.t55 IN_P.t1 bias21.t36 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X122 m9m10.t458 bias1.t108 VCC.t958 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X123 VCC.t957 bias1.t109 m1m2.t462 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X124 VCC.t956 bias1.t110 m1m2.t461 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X125 bias1.t6 VB_A.t7 m1m2.t516 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X126 m9m10.t457 bias1.t111 VCC.t955 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X127 a_46836_49340.t10 IN_P.t2 bias21.t35 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X128 a_46836_49340.t44 IN_M.t1 bias3.t29 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X129 dummy_3.t79 VB_B.t4 dummy_3.t78 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X130 m9m10.t456 bias1.t112 VCC.t954 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X131 VCC.t953 bias1.t113 m1m2.t460 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X132 VCC.t945 bias1.t114 m1m2.t459 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X133 dummy_9.t399 bias1.t115 dummy_9.t398 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X134 m9m10.t455 bias1.t116 VCC.t952 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X135 VCC.t951 bias1.t117 m1m2.t458 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X136 m9m10.t454 bias1.t118 VCC.t950 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X137 VCC.t949 bias1.t119 m1m2.t457 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X138 m9m10.t520 VB_A.t8 OUT.t27 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X139 m9m10.t453 bias1.t120 VCC.t948 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X140 VCC.t947 bias1.t121 m1m2.t456 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X141 VCC.t946 bias1.t122 m1m2.t455 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X142 VCC.t944 bias1.t123 m1m2.t454 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X143 bias1.t6 VB_A.t9 m1m2.t513 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X144 VCC.t943 bias1.t124 m1m2.t453 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X145 m11m12.t29 VB_B.t5 OUT.t48 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X146 m9m10.t452 bias1.t125 VCC.t942 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X147 dummy_2.t79 VB_A.t10 dummy_2.t78 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X148 m9m10.t451 bias1.t126 VCC.t941 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X149 VCC.t940 bias1.t127 m1m2.t452 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X150 dummy_9.t397 bias1.t128 dummy_9.t396 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X151 OUT.t59 VB_B.t6 m11m12.t28 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X152 m9m10.t450 bias1.t129 VCC.t939 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X153 VCC.t938 bias1.t130 m1m2.t451 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X154 dummy_9.t395 bias1.t131 dummy_9.t394 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X155 m9m10.t449 bias1.t132 VCC.t937 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X156 m9m10.t448 bias1.t133 VCC.t915 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X157 dummy_9.t393 bias1.t134 dummy_9.t392 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X158 VCC.t936 bias1.t135 m1m2.t450 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X159 m9m10.t447 bias1.t136 VCC.t935 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X160 VCC.t934 bias1.t137 m1m2.t449 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X161 m9m10.t446 bias1.t138 VCC.t933 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X162 dummy_3.t77 VB_B.t7 dummy_3.t76 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X163 VCC.t932 bias1.t139 m1m2.t448 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X164 bias21.t34 IN_P.t3 a_46836_49340.t11 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X165 m9m10.t518 VB_A.t11 OUT.t26 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X166 m9m10.t445 bias1.t140 VCC.t914 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X167 m9m10.t444 bias1.t141 VCC.t913 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X168 VCC.t931 bias1.t142 m1m2.t447 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X169 m9m10.t443 bias1.t143 VCC.t930 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X170 dummy_9.t391 bias1.t144 dummy_9.t390 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X171 dummy_9.t389 bias1.t145 dummy_9.t388 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X172 a_46836_49340.t62 IN_P.t4 bias21.t33 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X173 m9m10.t442 bias1.t146 VCC.t929 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X174 VCC.t928 bias1.t147 m1m2.t446 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X175 m9m10.t441 bias1.t148 VCC.t927 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X176 VCC.t926 bias1.t149 m1m2.t445 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X177 dummy_2.t77 VB_A.t12 dummy_2.t76 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X178 m9m10.t440 bias1.t150 VCC.t925 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X179 m9m10.t439 bias1.t151 VCC.t924 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X180 m9m10.t438 bias1.t152 VCC.t923 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X181 m9m10.t437 bias1.t153 VCC.t922 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X182 m9m10.t436 bias1.t154 VCC.t921 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X183 m9m10.t435 bias1.t155 VCC.t920 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X184 VCC.t919 bias1.t156 m1m2.t444 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X185 dummy_9.t387 bias1.t157 dummy_9.t386 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X186 OUT.t55 VB_B.t8 m11m12.t27 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X187 m9m10.t434 bias1.t158 VCC.t918 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X188 m9m10.t433 bias1.t159 VCC.t917 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X189 VCC.t916 bias1.t160 m1m2.t443 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X190 m9m10.t432 bias1.t161 VCC.t912 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X191 m9m10.t431 bias1.t162 VCC.t911 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X192 m9m10.t430 bias1.t163 VCC.t910 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X193 m9m10.t429 bias1.t164 VCC.t909 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X194 dummy_9.t385 bias1.t165 dummy_9.t384 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X195 m9m10.t428 bias1.t166 VCC.t908 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X196 VCC.t906 bias1.t167 m1m2.t442 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X197 VCC.t907 bias1.t168 m1m2.t441 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X198 dummy_9.t383 bias1.t169 dummy_9.t382 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X199 VCC.t905 bias1.t170 m1m2.t440 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X200 dummy_9.t381 bias1.t171 dummy_9.t380 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X201 m9m10.t427 bias1.t172 VCC.t904 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X202 dummy_4.t33 bias3.t41 dummy_4.t32 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X203 m9m10.t426 bias1.t173 VCC.t903 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X204 OUT.t25 VB_A.t13 m9m10.t517 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X205 m9m10.t425 bias1.t174 VCC.t902 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X206 dummy_9.t379 bias1.t175 dummy_9.t378 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X207 VCC.t901 bias1.t176 m1m2.t439 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X208 VCC.t900 bias1.t177 m1m2.t438 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X209 dummy_3.t75 VB_B.t9 dummy_3.t74 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X210 m9m10.t424 bias1.t178 VCC.t899 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X211 dummy_9.t377 bias1.t179 dummy_9.t376 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X212 m9m10.t423 bias1.t180 VCC.t898 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X213 VCC.t897 bias1.t181 m1m2.t437 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X214 m9m10.t422 bias1.t182 VCC.t896 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X215 VCC.t895 bias1.t183 m1m2.t436 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X216 m9m10.t421 bias1.t184 VCC.t894 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X217 dummy_9.t375 bias1.t185 dummy_9.t374 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X218 m9m10.t420 bias1.t186 VCC.t893 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X219 m9m10.t419 bias1.t187 VCC.t892 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X220 m9m10.t418 bias1.t188 VCC.t889 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X221 m9m10.t417 bias1.t189 VCC.t891 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X222 VCC.t890 bias1.t190 m1m2.t435 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X223 VCC.t888 bias1.t191 m1m2.t434 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X224 dummy_9.t373 bias1.t192 dummy_9.t372 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X225 dummy_2.t75 VB_A.t14 dummy_2.t74 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X226 m9m10.t416 bias1.t193 VCC.t887 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X227 m9m10.t415 bias1.t194 VCC.t886 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X228 OUT.t24 VB_A.t15 m9m10.t514 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X229 VCC.t885 bias1.t195 m1m2.t433 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X230 m9m10.t414 bias1.t196 VCC.t884 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X231 OUT.t56 VB_B.t10 m11m12.t26 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X232 dummy_9.t371 bias1.t197 dummy_9.t370 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X233 dummy_2.t73 VB_A.t16 dummy_2.t72 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X234 OUT.t54 VB_B.t11 m11m12.t25 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X235 m9m10.t413 bias1.t198 VCC.t883 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X236 m9m10.t412 bias1.t199 VCC.t882 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X237 VCC.t881 bias1.t200 m1m2.t432 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X238 m9m10.t411 bias1.t201 VCC.t880 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X239 VCC.t879 bias1.t202 m1m2.t431 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X240 VCC.t878 bias1.t203 m1m2.t430 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X241 VCC.t877 bias1.t204 m1m2.t429 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X242 m9m10.t410 bias1.t205 VCC.t876 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X243 VCC.t875 bias1.t206 m1m2.t428 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X244 dummy_9.t369 bias1.t207 dummy_9.t368 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X245 dummy_3.t73 VB_B.t12 dummy_3.t72 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X246 VCC.t874 bias1.t208 m1m2.t427 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X247 m9m10.t409 bias1.t209 VCC.t873 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X248 m9m10.t408 bias1.t210 VCC.t872 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X249 m9m10.t407 bias1.t211 VCC.t871 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X250 m9m10.t406 bias1.t212 VCC.t870 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X251 m9m10.t405 bias1.t213 VCC.t869 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X252 dummy_9.t367 bias1.t214 dummy_9.t366 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X253 m9m10.t404 bias1.t215 VCC.t868 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X254 VCC.t867 bias1.t216 m1m2.t426 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X255 m9m10.t403 bias1.t217 VCC.t863 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X256 m9m10.t402 bias1.t218 VCC.t866 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X257 VCC.t865 bias1.t219 m1m2.t425 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X258 m9m10.t401 bias1.t220 VCC.t864 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X259 VCC.t862 bias1.t221 m1m2.t424 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X260 VCC.t861 bias1.t222 m1m2.t423 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X261 a_46836_49340.t43 IN_M.t2 bias3.t12 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X262 VCC.t860 bias1.t223 m1m2.t422 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X263 m9m10.t400 bias1.t224 VCC.t859 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X264 m9m10.t399 bias1.t225 VCC.t858 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X265 a_46836_49340.t42 IN_M.t3 bias3.t13 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X266 VCC.t857 bias1.t226 m1m2.t421 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X267 m9m10.t398 bias1.t227 VCC.t855 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X268 VCC.t856 bias1.t228 m1m2.t420 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X269 m9m10.t397 bias1.t229 VCC.t854 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X270 VCC.t853 bias1.t230 m1m2.t419 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X271 dummy_9.t365 bias1.t231 dummy_9.t364 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X272 m11m12.t24 VB_B.t13 OUT.t58 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X273 VCC.t852 bias1.t232 m1m2.t418 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X274 dummy_9.t363 bias1.t233 dummy_9.t362 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X275 m9m10.t396 bias1.t234 VCC.t851 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X276 VCC.t850 bias1.t235 m1m2.t417 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X277 dummy_9.t361 bias1.t236 dummy_9.t360 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X278 m9m10.t395 bias1.t237 VCC.t849 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X279 m9m10.t394 bias1.t238 VCC.t848 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X280 m9m10.t393 bias1.t239 VCC.t847 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X281 VCC.t846 bias1.t240 m1m2.t416 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X282 VCC.t786 bias1.t241 m1m2.t415 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X283 VCC.t845 bias1.t242 m1m2.t414 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X284 m9m10.t392 bias1.t243 VCC.t844 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X285 VCC.t843 bias1.t244 m1m2.t413 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X286 VCC.t842 bias1.t245 m1m2.t412 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X287 m9m10.t391 bias1.t246 VCC.t841 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X288 VCC.t840 bias1.t247 m1m2.t411 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X289 dummy_100.t33 IB.t11 dummy_100.t32 VCC.t1038 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X290 m9m10.t515 VB_A.t17 OUT.t23 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X291 a_46836_49340.t41 IN_M.t4 bias3.t20 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X292 dummy_3.t71 VB_B.t14 dummy_3.t70 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X293 m9m10.t390 bias1.t248 VCC.t839 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X294 dummy_9.t359 bias1.t249 dummy_9.t358 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X295 bias1.t6 VB_A.t18 m1m2.t509 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X296 m9m10.t389 bias1.t250 VCC.t838 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X297 VCC.t837 bias1.t251 m1m2.t410 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X298 m9m10.t388 bias1.t252 VCC.t836 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X299 dummy_9.t357 bias1.t253 dummy_9.t356 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X300 dummy_9.t355 bias1.t254 dummy_9.t354 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X301 m9m10.t387 bias1.t255 VCC.t832 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X302 dummy_3.t69 VB_B.t15 dummy_3.t68 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X303 m9m10.t386 bias1.t256 VCC.t835 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X304 VCC.t834 bias1.t257 m1m2.t409 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X305 VCC.t833 bias1.t258 m1m2.t408 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X306 m9m10.t385 bias1.t259 VCC.t831 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X307 VCC.t830 bias1.t260 m1m2.t407 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X308 m9m10.t384 bias1.t261 VCC.t829 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X309 VCC.t828 bias1.t262 m1m2.t406 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X310 m9m10.t383 bias1.t263 VCC.t827 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X311 dummy_9.t353 bias1.t207 dummy_9.t352 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X312 bias3.t21 IN_M.t5 a_46836_49340.t40 VCC.t9 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X313 VCC.t826 bias1.t264 m1m2.t405 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X314 dummy_9.t351 bias1.t265 dummy_9.t350 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X315 VCC.t825 bias1.t266 m1m2.t404 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X316 dummy_9.t349 bias1.t267 dummy_9.t348 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X317 m9m10.t382 bias1.t268 VCC.t824 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X318 dummy_9.t347 bias1.t269 dummy_9.t346 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X319 VCC.t823 bias1.t270 m1m2.t403 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X320 m9m10.t381 bias1.t271 VCC.t822 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X321 m9m10.t380 bias1.t272 VCC.t816 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X322 VCC.t821 bias1.t273 m1m2.t402 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X323 m1m2.t510 VB_A.t19 bias1.t6 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X324 m9m10.t379 bias1.t274 VCC.t820 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X325 dummy_3.t67 VB_B.t16 dummy_3.t66 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X326 m9m10.t378 bias1.t275 VCC.t819 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X327 VCC.t818 bias1.t276 m1m2.t401 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X328 OUT.t52 VB_B.t17 m11m12.t23 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X329 m9m10.t377 bias1.t277 VCC.t817 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X330 m9m10.t376 bias1.t278 VCC.t815 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X331 dummy_2.t71 VB_A.t20 dummy_2.t70 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X332 m9m10.t375 bias1.t279 VCC.t814 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X333 dummy_100.t31 IB.t12 dummy_100.t30 VCC.t2 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X334 dummy_2.t69 VB_A.t21 dummy_2.t68 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X335 dummy_9.t345 bias1.t280 dummy_9.t344 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X336 dummy_9.t343 bias1.t281 dummy_9.t342 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X337 bias3.t34 IN_M.t6 a_46836_49340.t39 VCC.t9 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X338 VCC.t813 bias1.t282 m1m2.t400 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X339 dummy_9.t341 bias1.t283 dummy_9.t340 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X340 m9m10.t374 bias1.t284 VCC.t812 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X341 dummy_3.t65 VB_B.t18 dummy_3.t64 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X342 VCC.t811 bias1.t285 m1m2.t399 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X343 m9m10.t373 bias1.t286 VCC.t810 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X344 VSS.t13 bias3.t42 m3m4.t30 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=1
**devattr s=58000,2116 d=58000,2116
X345 VCC.t809 bias1.t287 m1m2.t398 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X346 m9m10.t372 bias1.t288 VCC.t808 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X347 VCC.t805 bias1.t289 m1m2.t397 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X348 m9m10.t371 bias1.t290 VCC.t807 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X349 dummy_3.t63 VB_B.t19 dummy_3.t62 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X350 VCC.t806 bias1.t291 m1m2.t396 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X351 m9m10.t511 VB_A.t22 OUT.t22 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X352 m9m10.t370 bias1.t292 VCC.t804 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X353 dummy_9.t339 bias1.t293 dummy_9.t338 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X354 VCC.t803 bias1.t294 m1m2.t395 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X355 VCC.t802 bias1.t295 m1m2.t394 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X356 dummy_9.t337 bias1.t296 dummy_9.t336 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X357 dummy_9.t335 bias1.t297 dummy_9.t334 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X358 VCC.t787 bias1.t298 m1m2.t393 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X359 m9m10.t369 bias1.t299 VCC.t801 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X360 m9m10.t368 bias1.t300 VCC.t800 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X361 m11m12.t22 VB_B.t20 OUT.t39 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X362 VCC.t799 bias1.t301 m1m2.t392 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X363 m9m10.t367 bias1.t302 VCC.t798 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X364 dummy_9.t333 bias1.t303 dummy_9.t332 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X365 dummy_2.t67 VB_A.t23 dummy_2.t66 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X366 bias3.t35 IN_M.t7 a_46836_49340.t38 VCC.t9 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X367 m9m10.t366 bias1.t304 VCC.t797 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X368 m9m10.t365 bias1.t305 VCC.t796 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X369 dummy_9.t331 bias1.t306 dummy_9.t330 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X370 m9m10.t364 bias1.t307 VCC.t795 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X371 VCC.t794 bias1.t308 m1m2.t391 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X372 VCC.t793 bias1.t309 m1m2.t390 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X373 VCC.t792 bias1.t310 m1m2.t389 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X374 dummy_9.t329 bias1.t311 dummy_9.t328 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X375 m9m10.t363 bias1.t312 VCC.t791 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X376 dummy_9.t327 bias1.t313 dummy_9.t326 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X377 m9m10.t362 bias1.t314 VCC.t790 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X378 dummy_3.t61 VB_B.t21 dummy_3.t60 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X379 VCC.t789 bias1.t315 m1m2.t388 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X380 m9m10.t361 bias1.t316 VCC.t788 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X381 VCC.t785 bias1.t317 m1m2.t387 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X382 dummy_3.t59 VB_B.t22 dummy_3.t58 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X383 m9m10.t360 bias1.t318 VCC.t784 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X384 dummy_9.t325 bias1.t319 dummy_9.t324 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X385 dummy_9.t323 bias1.t320 dummy_9.t322 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X386 dummy_2.t65 VB_A.t24 dummy_2.t64 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X387 dummy_9.t321 bias1.t321 dummy_9.t320 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X388 dummy_9.t319 bias1.t57 dummy_9.t318 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X389 m9m10.t359 bias1.t322 VCC.t783 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X390 m9m10.t358 bias1.t323 VCC.t782 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X391 m9m10.t357 bias1.t324 VCC.t781 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X392 dummy_4.t31 bias3.t43 dummy_4.t30 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X393 m9m10.t356 bias1.t325 VCC.t780 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X394 VCC.t779 bias1.t326 m1m2.t386 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X395 dummy_9.t317 bias1.t327 dummy_9.t316 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X396 VCC.t773 bias1.t328 m1m2.t385 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X397 VCC.t778 bias1.t329 m1m2.t384 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X398 m9m10.t355 bias1.t330 VCC.t777 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X399 VCC.t776 bias1.t331 m1m2.t383 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X400 m9m10.t354 bias1.t332 VCC.t775 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X401 dummy_9.t315 bias1.t333 dummy_9.t314 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X402 VCC.t774 bias1.t334 m1m2.t382 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X403 m9m10.t353 bias1.t335 VCC.t772 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X404 VCC.t771 bias1.t336 m1m2.t381 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X405 dummy_100.t29 IB.t13 dummy_100.t28 VCC.t8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X406 dummy_3.t57 VB_B.t23 dummy_3.t56 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X407 VCC.t770 bias1.t337 m1m2.t380 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X408 dummy_9.t313 bias1.t338 dummy_9.t312 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X409 m9m10.t352 bias1.t339 VCC.t769 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X410 m9m10.t351 bias1.t340 VCC.t768 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X411 VCC.t767 bias1.t341 m1m2.t379 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X412 OUT.t31 VB_B.t24 m11m12.t21 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X413 VCC.t766 bias1.t342 m1m2.t378 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X414 VCC.t764 bias1.t343 m1m2.t377 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X415 dummy_9.t311 bias1.t344 dummy_9.t310 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X416 dummy_2.t63 VB_A.t25 dummy_2.t62 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X417 m9m10.t350 bias1.t345 VCC.t765 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X418 m9m10.t349 bias1.t346 VCC.t763 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X419 VCC.t762 bias1.t347 m1m2.t376 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X420 VCC.t761 bias1.t348 m1m2.t375 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X421 bias1.t5 VB_B.t25 m3m4.t27 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X422 m9m10.t348 bias1.t349 VCC.t760 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X423 m9m10.t347 bias1.t350 VCC.t759 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X424 VCC.t758 bias1.t351 m1m2.t374 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X425 m9m10.t509 VB_A.t26 OUT.t21 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X426 m9m10.t346 bias1.t352 VCC.t743 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X427 m9m10.t345 bias1.t353 VCC.t757 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X428 VCC.t756 bias1.t354 m1m2.t373 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X429 m9m10.t344 bias1.t355 VCC.t755 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X430 dummy_100.t27 IB.t14 dummy_100.t26 VCC.t8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X431 VCC.t754 bias1.t356 m1m2.t372 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X432 m9m10.t343 bias1.t357 VCC.t753 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X433 bias3.t36 IN_M.t8 a_46836_49340.t37 VCC.t9 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X434 m9m10.t342 bias1.t358 VCC.t752 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X435 dummy_9.t309 bias1.t359 dummy_9.t308 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X436 VCC.t751 bias1.t360 m1m2.t371 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X437 m9m10.t341 bias1.t361 VCC.t739 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X438 m9m10.t340 bias1.t362 VCC.t750 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X439 m9m10.t339 bias1.t363 VCC.t749 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X440 VCC.t748 bias1.t364 m1m2.t370 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X441 a_46836_49340.t36 IN_M.t9 bias3.t37 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X442 VCC.t741 bias1.t365 m1m2.t369 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X443 VCC.t747 bias1.t366 m1m2.t368 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X444 a_46836_49340.t35 IN_M.t10 bias3.t14 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X445 VCC.t740 bias1.t367 m1m2.t367 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X446 VCC.t746 bias1.t368 m1m2.t366 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X447 dummy_9.t307 bias1.t369 dummy_9.t306 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X448 VCC.t745 bias1.t370 m1m2.t365 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X449 VCC.t744 bias1.t371 m1m2.t364 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X450 dummy_9.t305 bias1.t372 dummy_9.t304 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X451 VCC.t742 bias1.t373 m1m2.t363 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X452 dummy_9.t303 bias1.t374 dummy_9.t302 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X453 VCC.t738 bias1.t375 m1m2.t362 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X454 m9m10.t338 bias1.t376 VCC.t737 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X455 VCC.t736 bias1.t377 m1m2.t361 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X456 dummy_9.t301 bias1.t378 dummy_9.t300 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X457 m9m10.t337 bias1.t379 VCC.t735 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X458 VCC.t734 bias1.t380 m1m2.t360 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X459 VCC.t731 bias1.t381 m1m2.t359 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X460 VCC.t733 bias1.t382 m1m2.t358 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X461 VCC.t732 bias1.t383 m1m2.t357 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X462 m9m10.t336 bias1.t384 VCC.t730 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X463 bias1.t6 VB_A.t27 m1m2.t506 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X464 a_46836_49340.t63 IN_P.t5 bias21.t32 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X465 dummy_2.t61 VB_A.t28 dummy_2.t60 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X466 dummy_3.t55 VB_B.t26 dummy_3.t54 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X467 VCC.t729 bias1.t385 m1m2.t356 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X468 VCC.t728 bias1.t386 m1m2.t355 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X469 m9m10.t335 bias1.t387 VCC.t727 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X470 dummy_9.t299 bias1.t388 dummy_9.t298 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X471 m9m10.t334 bias1.t389 VCC.t726 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X472 m9m10.t333 bias1.t390 VCC.t725 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X473 VCC.t724 bias1.t391 m1m2.t354 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X474 VSS.t17 bias3.t6 bias3.t7 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X475 VCC.t675 bias1.t392 m1m2.t353 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X476 bias21.t31 IN_P.t6 a_46836_49340.t58 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X477 m9m10.t506 VB_A.t29 OUT.t20 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X478 m9m10.t332 bias1.t393 VCC.t676 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X479 VCC.t723 bias1.t394 m1m2.t352 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X480 VCC.t722 bias1.t395 m1m2.t351 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X481 m9m10.t331 bias1.t396 VCC.t721 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X482 dummy_9.t297 bias1.t397 dummy_9.t296 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X483 bias3.t15 IN_M.t11 a_46836_49340.t34 VCC.t9 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X484 m9m10.t330 bias1.t398 VCC.t720 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X485 VCC.t719 bias1.t399 m1m2.t350 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X486 dummy_2.t59 VB_A.t30 dummy_2.t58 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X487 VCC.t718 bias1.t400 m1m2.t349 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X488 VSS.t18 bias3.t4 bias3.t5 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X489 dummy_9.t295 bias1.t401 dummy_9.t294 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X490 dummy_3.t53 VB_B.t27 dummy_3.t52 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X491 VCC.t717 bias1.t402 m1m2.t348 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X492 VCC.t716 bias1.t403 m1m2.t347 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X493 dummy_4.t29 bias3.t44 dummy_4.t28 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X494 m9m10.t329 bias1.t404 VCC.t715 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X495 m9m10.t328 bias1.t405 VCC.t714 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X496 VCC.t713 bias1.t406 m1m2.t346 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X497 bias1.t6 VB_A.t31 m1m2.t505 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X498 VCC.t710 bias1.t407 m1m2.t345 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X499 m9m10.t327 bias1.t408 VCC.t712 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X500 VCC.t711 bias1.t409 m1m2.t344 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X501 a_46836_49340.t33 IN_M.t12 bias3.t16 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X502 OUT.t19 VB_A.t32 m9m10.t504 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X503 dummy_4.t27 bias3.t45 dummy_4.t26 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X504 m9m10.t326 bias1.t410 VCC.t709 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X505 VCC.t708 bias1.t411 m1m2.t343 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X506 VCC.t707 bias1.t412 m1m2.t342 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X507 bias21.t30 IN_P.t7 a_46836_49340.t59 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X508 m9m10.t325 bias1.t413 VCC.t706 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X509 m9m10.t324 bias1.t414 VCC.t705 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X510 VCC.t703 bias1.t415 m1m2.t341 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X511 dummy_9.t293 bias1.t416 dummy_9.t292 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X512 m3m4.t26 VB_B.t28 bias1.t4 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X513 dummy_9.t291 bias1.t417 dummy_9.t290 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X514 VCC.t704 bias1.t418 m1m2.t340 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X515 m9m10.t323 bias1.t419 VCC.t702 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X516 VCC.t10 IB.t15 a_46836_49340.t51 VCC.t2 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X517 a_46836_49340.t50 IB.t16 VCC.t1 VCC.t0 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X518 m9m10.t322 bias1.t420 VCC.t701 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X519 VCC.t700 bias1.t421 m1m2.t339 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X520 m9m10.t321 bias1.t422 VCC.t699 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X521 VCC.t3 IB.t17 a_46836_49340.t49 VCC.t2 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X522 VCC.t698 bias1.t423 m1m2.t338 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X523 bias1.t6 VB_A.t33 m1m2.t501 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X524 dummy_9.t289 bias1.t424 dummy_9.t288 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X525 m9m10.t320 bias1.t425 VCC.t697 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X526 dummy_3.t51 VB_B.t29 dummy_3.t50 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X527 m11m12.t20 VB_B.t30 OUT.t40 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X528 dummy_3.t49 VB_B.t31 dummy_3.t48 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X529 dummy_9.t287 bias1.t426 dummy_9.t286 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X530 m9m10.t319 bias1.t427 VCC.t696 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X531 m9m10.t318 bias1.t428 VCC.t695 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X532 m9m10.t317 bias1.t429 VCC.t694 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X533 m9m10.t316 bias1.t430 VCC.t691 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X534 dummy_9.t285 bias1.t431 dummy_9.t284 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X535 m9m10.t315 bias1.t432 VCC.t690 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X536 VCC.t693 bias1.t433 m1m2.t337 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X537 dummy_100.t25 IB.t18 dummy_100.t24 VCC.t2 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X538 dummy_9.t283 bias1.t434 dummy_9.t282 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X539 m9m10.t314 bias1.t435 VCC.t692 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X540 VCC.t689 bias1.t436 m1m2.t336 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X541 dummy_4.t25 bias3.t46 dummy_4.t24 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X542 m9m10.t313 bias1.t437 VCC.t688 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X543 VCC.t687 bias1.t438 m1m2.t335 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X544 bias21.t29 IN_P.t8 a_46836_49340.t2 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X545 m9m10.t312 bias1.t439 VCC.t686 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X546 dummy_3.t47 VB_B.t32 dummy_3.t46 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X547 VCC.t685 bias1.t440 m1m2.t334 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X548 dummy_9.t281 bias1.t441 dummy_9.t280 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X549 m9m10.t311 bias1.t442 VCC.t684 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X550 m9m10.t310 bias1.t443 VCC.t683 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X551 m9m10.t309 bias1.t444 VCC.t682 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X552 dummy_9.t279 bias1.t445 dummy_9.t278 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X553 m9m10.t308 bias1.t446 VCC.t681 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X554 m3m4.t25 VB_B.t33 bias1.t1 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X555 dummy_9.t277 bias1.t447 dummy_9.t276 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X556 m1m2.t502 VB_A.t34 bias1.t6 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X557 VCC.t680 bias1.t448 m1m2.t333 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X558 VCC.t679 bias1.t449 m1m2.t332 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X559 dummy_9.t275 bias1.t450 dummy_9.t274 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X560 m9m10.t307 bias1.t451 VCC.t678 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X561 dummy_3.t45 VB_B.t34 dummy_3.t44 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X562 VSS.t16 bias3.t2 bias3.t3 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X563 m9m10.t306 bias1.t452 VCC.t677 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X564 m9m10.t305 bias1.t453 VCC.t674 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X565 VCC.t673 bias1.t454 m1m2.t331 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X566 dummy_9.t273 bias1.t455 dummy_9.t272 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X567 m9m10.t304 bias1.t456 VCC.t672 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X568 VCC.t670 bias1.t457 m1m2.t330 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X569 m9m10.t303 bias1.t458 VCC.t671 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X570 m9m10.t302 bias1.t459 VCC.t669 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X571 m9m10.t301 bias1.t460 VCC.t668 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X572 dummy_9.t271 bias1.t461 dummy_9.t270 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X573 m11m12.t19 VB_B.t35 OUT.t49 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X574 VCC.t667 bias1.t462 m1m2.t329 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X575 dummy_2.t57 VB_A.t35 dummy_2.t56 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X576 m9m10.t300 bias1.t463 VCC.t666 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X577 dummy_9.t269 bias1.t231 dummy_9.t268 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X578 VCC.t665 bias1.t464 m1m2.t328 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X579 m9m10.t299 bias1.t465 VCC.t664 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X580 dummy_9.t267 bias1.t231 dummy_9.t266 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X581 m9m10.t298 bias1.t466 VCC.t544 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X582 m9m10.t297 bias1.t467 VCC.t663 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X583 dummy_3.t43 VB_B.t36 dummy_3.t42 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X584 m9m10.t296 bias1.t468 VCC.t662 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X585 m9m10.t295 bias1.t469 VCC.t661 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X586 dummy_9.t265 bias1.t470 dummy_9.t264 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X587 VCC.t660 bias1.t471 m1m2.t327 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X588 dummy_9.t263 bias1.t472 dummy_9.t262 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X589 VCC.t659 bias1.t473 m1m2.t326 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X590 OUT.t41 VB_B.t37 m11m12.t18 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X591 m9m10.t294 bias1.t474 VCC.t658 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X592 VCC.t657 bias1.t475 m1m2.t325 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X593 dummy_9.t261 bias1.t476 dummy_9.t260 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X594 dummy_100.t23 IB.t19 dummy_100.t22 VCC.t7 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X595 dummy_9.t259 bias1.t477 dummy_9.t258 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X596 dummy_3.t41 VB_B.t38 dummy_3.t40 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X597 VCC.t656 bias1.t478 m1m2.t324 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X598 VCC.t655 bias1.t479 m1m2.t323 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X599 m9m10.t293 bias1.t480 VCC.t654 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X600 m9m10.t292 bias1.t481 VCC.t650 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X601 VCC.t653 bias1.t482 m1m2.t322 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X602 VCC.t652 bias1.t483 m1m2.t321 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X603 dummy_3.t39 VB_B.t39 dummy_3.t38 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X604 dummy_9.t257 bias1.t484 dummy_9.t256 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X605 VCC.t651 bias1.t485 m1m2.t320 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X606 dummy_9.t255 bias1.t486 dummy_9.t254 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X607 VCC.t649 bias1.t487 m1m2.t319 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X608 dummy_9.t253 bias1.t231 dummy_9.t252 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X609 m9m10.t291 bias1.t488 VCC.t648 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X610 VCC.t647 bias1.t489 m1m2.t318 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X611 dummy_9.t251 bias1.t490 dummy_9.t250 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X612 dummy_9.t249 bias1.t491 dummy_9.t248 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X613 m3m4.t24 VB_B.t40 bias1.t4 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X614 dummy_2.t55 VB_A.t36 dummy_2.t54 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X615 m3m4.t23 VB_B.t41 bias1.t5 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X616 m9m10.t290 bias1.t492 VCC.t646 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X617 VCC.t645 bias1.t493 m1m2.t317 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X618 m9m10.t289 bias1.t494 VCC.t644 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X619 m9m10.t288 bias1.t495 VCC.t643 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X620 VCC.t642 bias1.t496 m1m2.t316 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X621 VCC.t635 bias1.t497 m1m2.t315 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X622 VCC.t641 bias1.t498 m1m2.t314 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X623 bias21.t28 IN_P.t9 a_46836_49340.t3 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X624 dummy_4.t23 bias3.t47 dummy_4.t22 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X625 m9m10.t287 bias1.t499 VCC.t640 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X626 dummy_9.t247 bias1.t500 dummy_9.t246 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X627 dummy_2.t53 VB_A.t37 dummy_2.t52 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X628 VCC.t639 bias1.t501 m1m2.t313 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X629 m9m10.t286 bias1.t502 VCC.t638 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X630 m11m12.t17 VB_B.t42 OUT.t51 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X631 dummy_3.t37 VB_B.t43 dummy_3.t36 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X632 VCC.t636 bias1.t503 m1m2.t312 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X633 m9m10.t285 bias1.t504 VCC.t637 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X634 m9m10.t284 bias1.t505 VCC.t634 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X635 dummy_9.t245 bias1.t506 dummy_9.t244 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X636 dummy_9.t243 bias1.t507 dummy_9.t242 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X637 VCC.t633 bias1.t508 m1m2.t311 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X638 VCC.t632 bias1.t509 m1m2.t310 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X639 m9m10.t283 bias1.t510 VCC.t631 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X640 m9m10.t282 bias1.t511 VCC.t630 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X641 m9m10.t281 bias1.t512 VCC.t629 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X642 VCC.t628 bias1.t513 m1m2.t309 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X643 VCC.t627 bias1.t514 m1m2.t308 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X644 m9m10.t280 bias1.t515 VCC.t626 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X645 bias3.t17 IN_M.t13 a_46836_49340.t32 VCC.t9 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X646 VCC.t622 bias1.t516 m1m2.t307 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X647 dummy_3.t35 VB_B.t44 dummy_3.t34 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X648 bias3.t18 IN_M.t14 a_46836_49340.t31 VCC.t9 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X649 dummy_100.t21 IB.t20 dummy_100.t20 VCC.t6 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X650 dummy_9.t241 bias1.t517 dummy_9.t240 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X651 dummy_9.t239 bias1.t518 dummy_9.t238 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X652 OUT.t30 VB_B.t45 m11m12.t16 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X653 m9m10.t279 bias1.t519 VCC.t625 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X654 VCC.t624 bias1.t520 m1m2.t306 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X655 VCC.t621 bias1.t521 m1m2.t305 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X656 m9m10.t278 bias1.t522 VCC.t623 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X657 m9m10.t529 VB_A.t38 OUT.t18 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X658 m9m10.t277 bias1.t523 VCC.t620 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X659 VCC.t619 bias1.t524 m1m2.t304 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X660 VCC.t607 bias1.t525 m1m2.t303 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X661 VCC.t618 bias1.t526 m1m2.t302 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X662 VCC.t617 bias1.t527 m1m2.t301 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X663 VCC.t616 bias1.t528 m1m2.t300 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X664 bias1.t6 VB_A.t39 m1m2.t529 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X665 dummy_4.t21 bias3.t48 dummy_4.t20 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X666 VCC.t615 bias1.t529 m1m2.t299 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X667 bias3.t19 IN_M.t15 a_46836_49340.t30 VCC.t9 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X668 m9m10.t276 bias1.t530 VCC.t614 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X669 m9m10.t275 bias1.t531 VCC.t613 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X670 dummy_9.t237 bias1.t532 dummy_9.t236 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X671 VCC.t612 bias1.t533 m1m2.t298 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X672 VCC.t606 bias1.t534 m1m2.t297 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X673 dummy_3.t33 VB_B.t46 dummy_3.t32 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X674 VCC.t611 bias1.t535 m1m2.t296 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X675 VCC.t610 bias1.t536 m1m2.t295 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X676 bias21.t27 IN_P.t10 a_46836_49340.t56 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X677 m9m10.t528 VB_A.t40 OUT.t17 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X678 m9m10.t274 bias1.t537 VCC.t609 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X679 m9m10.t273 bias1.t538 VCC.t608 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X680 m9m10.t272 bias1.t539 VCC.t605 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X681 m9m10.t271 bias1.t540 VCC.t604 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X682 m9m10.t270 bias1.t541 VCC.t603 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X683 m9m10.t269 bias1.t542 VCC.t602 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X684 VCC.t601 bias1.t543 m1m2.t294 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X685 VCC.t598 bias1.t544 m1m2.t293 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X686 m9m10.t268 bias1.t545 VCC.t600 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X687 VCC.t599 bias1.t546 m1m2.t292 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X688 m9m10.t267 bias1.t547 VCC.t597 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X689 m9m10.t266 bias1.t548 VCC.t596 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X690 VCC.t595 bias1.t549 m1m2.t291 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X691 dummy_2.t51 VB_A.t41 dummy_2.t50 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X692 VCC.t594 bias1.t550 m1m2.t290 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X693 m3m4.t22 VB_B.t47 bias1.t3 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X694 dummy_9.t235 bias1.t551 dummy_9.t234 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X695 m9m10.t265 bias1.t552 VCC.t593 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X696 VCC.t592 bias1.t553 m1m2.t289 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X697 dummy_9.t233 bias1.t554 dummy_9.t232 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X698 dummy_9.t231 bias1.t555 dummy_9.t230 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X699 m9m10.t264 bias1.t556 VCC.t591 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X700 m9m10.t263 bias1.t557 VCC.t590 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X701 VCC.t586 bias1.t558 m1m2.t288 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X702 m9m10.t262 bias1.t559 VCC.t589 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X703 VCC.t588 bias1.t560 m1m2.t287 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X704 m9m10.t261 bias1.t561 VCC.t587 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X705 m9m10.t260 bias1.t562 VCC.t585 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X706 a_46836_49340.t57 IN_P.t11 bias21.t26 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X707 m11m12.t15 VB_B.t48 OUT.t44 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X708 VCC.t584 bias1.t563 m1m2.t286 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X709 bias1.t6 VB_A.t42 m1m2.t527 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X710 dummy_9.t229 bias1.t564 dummy_9.t228 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X711 dummy_2.t49 VB_A.t43 dummy_2.t48 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X712 m9m10.t259 bias1.t565 VCC.t583 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X713 VCC.t582 bias1.t566 m1m2.t285 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X714 m9m10.t258 bias1.t567 VCC.t581 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X715 m9m10.t257 bias1.t568 VCC.t580 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X716 m9m10.t256 bias1.t569 VCC.t579 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X717 VCC.t578 bias1.t570 m1m2.t284 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X718 dummy_9.t227 bias1.t571 dummy_9.t226 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X719 dummy_3.t31 VB_B.t49 dummy_3.t30 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X720 m9m10.t255 bias1.t572 VCC.t577 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X721 VCC.t574 bias1.t573 m1m2.t283 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X722 VCC.t576 bias1.t574 m1m2.t282 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X723 m9m10.t254 bias1.t575 VCC.t575 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X724 m9m10.t253 bias1.t576 VCC.t573 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X725 VCC.t572 bias1.t577 m1m2.t281 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X726 m1m2.t528 VB_A.t44 bias1.t6 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X727 VCC.t571 bias1.t578 m1m2.t280 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X728 dummy_9.t225 bias1.t579 dummy_9.t224 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X729 OUT.t32 VB_B.t50 m11m12.t14 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X730 VCC.t570 bias1.t580 m1m2.t279 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X731 VCC.t546 bias1.t581 m1m2.t278 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X732 m9m10.t252 bias1.t582 VCC.t569 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X733 dummy_9.t223 bias1.t583 dummy_9.t222 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X734 dummy_9.t221 bias1.t584 dummy_9.t220 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X735 m9m10.t251 bias1.t585 VCC.t568 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X736 VCC.t567 bias1.t586 m1m2.t277 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X737 dummy_9.t219 bias1.t587 dummy_9.t218 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X738 OUT.t16 VB_A.t45 m9m10.t527 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X739 m1m2.t525 VB_A.t46 bias1.t6 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X740 m9m10.t250 bias1.t588 VCC.t566 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X741 m9m10.t249 bias1.t589 VCC.t565 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X742 m9m10.t248 bias1.t590 VCC.t564 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X743 VCC.t545 bias1.t591 m1m2.t276 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X744 m9m10.t247 bias1.t592 VCC.t563 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X745 dummy_9.t217 bias1.t593 dummy_9.t216 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X746 dummy_3.t29 VB_B.t51 dummy_3.t28 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X747 VCC.t561 bias1.t594 m1m2.t275 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X748 VCC.t562 bias1.t595 m1m2.t274 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X749 VCC.t560 bias1.t596 m1m2.t273 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X750 dummy_9.t215 bias1.t207 dummy_9.t214 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X751 VCC.t559 bias1.t597 m1m2.t272 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X752 VCC.t558 bias1.t598 m1m2.t271 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X753 dummy_9.t213 bias1.t207 dummy_9.t212 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X754 VCC.t547 bias1.t599 m1m2.t270 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X755 m9m10.t246 bias1.t600 VCC.t557 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X756 VCC.t556 bias1.t601 m1m2.t269 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X757 m9m10.t245 bias1.t602 VCC.t555 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X758 dummy_9.t211 bias1.t603 dummy_9.t210 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X759 m1m2.t526 VB_A.t47 bias1.t6 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X760 dummy_2.t47 VB_A.t48 dummy_2.t46 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X761 VCC.t554 bias1.t604 m1m2.t268 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X762 dummy_9.t209 bias1.t605 dummy_9.t208 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X763 VCC.t553 bias1.t606 m1m2.t267 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X764 dummy_9.t207 bias1.t607 dummy_9.t206 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X765 VCC.t552 bias1.t608 m1m2.t266 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X766 VCC.t551 bias1.t609 m1m2.t265 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X767 VCC.t548 bias1.t610 m1m2.t264 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X768 m9m10.t244 bias1.t611 VCC.t550 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X769 dummy_9.t205 bias1.t612 dummy_9.t204 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X770 IB.t7 IB.t6 VCC.t1047 VCC.t7 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X771 VCC.t549 bias1.t613 m1m2.t263 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X772 VCC.t543 bias1.t614 m1m2.t262 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X773 m9m10.t243 bias1.t615 VCC.t542 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X774 IB.t5 IB.t4 VCC.t12 VCC.t7 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X775 m3m4.t21 VB_B.t52 bias1.t3 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X776 VCC.t541 bias1.t616 m1m2.t261 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X777 VCC.t540 bias1.t617 m1m2.t260 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X778 m9m10.t242 bias1.t618 VCC.t539 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X779 VCC.t538 bias1.t619 m1m2.t259 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X780 dummy_9.t203 bias1.t620 dummy_9.t202 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X781 m9m10.t241 bias1.t621 VCC.t537 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X782 m9m10.t240 bias1.t622 VCC.t536 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X783 VCC.t535 bias1.t623 m1m2.t258 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X784 m9m10.t239 bias1.t624 VCC.t534 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X785 VCC.t533 bias1.t625 m1m2.t257 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X786 bias1.t6 VB_A.t49 m1m2.t524 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X787 dummy_9.t201 bias1.t626 dummy_9.t200 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X788 a_46836_49340.t29 IN_M.t16 bias3.t32 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X789 dummy_2.t45 VB_A.t50 dummy_2.t44 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X790 m9m10.t238 bias1.t627 VCC.t532 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X791 VCC.t531 bias1.t628 m1m2.t256 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X792 VCC.t530 bias1.t629 m1m2.t255 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X793 m9m10.t237 bias1.t630 VCC.t529 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X794 dummy_9.t199 bias1.t631 dummy_9.t198 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X795 VCC.t527 bias1.t632 m1m2.t254 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X796 VCC.t528 bias1.t633 m1m2.t253 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X797 bias21.t25 IN_P.t12 a_46836_49340.t6 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X798 VCC.t526 bias1.t634 m1m2.t252 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X799 m9m10.t236 bias1.t635 VCC.t525 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X800 VCC.t518 bias1.t636 m1m2.t251 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X801 bias21.t24 IN_P.t13 a_46836_49340.t7 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X802 m9m10.t235 bias1.t637 VCC.t524 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X803 dummy_100.t19 IB.t21 dummy_100.t18 VCC.t0 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X804 bias21.t7 bias21.t6 VSS.t21 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X805 dummy_9.t197 bias1.t638 dummy_9.t196 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X806 VCC.t523 bias1.t639 m1m2.t250 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X807 VCC.t522 bias1.t640 m1m2.t249 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X808 bias3.t33 IN_M.t17 a_46836_49340.t28 VCC.t9 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X809 bias3.t8 IN_M.t18 a_46836_49340.t27 VCC.t9 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X810 m9m10.t234 bias1.t641 VCC.t521 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X811 dummy_2.t43 VB_A.t51 dummy_2.t42 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X812 dummy_9.t195 bias1.t642 dummy_9.t194 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X813 dummy_9.t193 bias1.t643 dummy_9.t192 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X814 VCC.t520 bias1.t644 m1m2.t248 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X815 bias1.t5 VB_B.t53 m3m4.t20 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X816 bias21.t5 bias21.t4 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X817 dummy_9.t191 bias1.t645 dummy_9.t190 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X818 m9m10.t233 bias1.t646 VCC.t519 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X819 VCC.t517 bias1.t647 m1m2.t247 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X820 a_46836_49340.t0 IN_P.t14 bias21.t23 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X821 VCC.t516 bias1.t648 m1m2.t246 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X822 VCC.t515 bias1.t649 m1m2.t245 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X823 VCC.t514 bias1.t650 m1m2.t244 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X824 m9m10.t232 bias1.t651 VCC.t513 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X825 bias21.t22 IN_P.t15 a_46836_49340.t1 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X826 m9m10.t231 bias1.t652 VCC.t512 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X827 dummy_9.t189 bias1.t653 dummy_9.t188 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X828 dummy_9.t187 bias1.t654 dummy_9.t186 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X829 dummy_100.t17 IB.t22 dummy_100.t16 VCC.t1038 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X830 VCC.t511 bias1.t655 m1m2.t243 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X831 m9m10.t230 bias1.t656 VCC.t510 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X832 m9m10.t229 bias1.t657 VCC.t509 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X833 m9m10.t228 bias1.t658 VCC.t508 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X834 m9m10.t227 bias1.t659 VCC.t499 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X835 VCC.t507 bias1.t660 m1m2.t242 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X836 VCC.t506 bias1.t661 m1m2.t241 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X837 bias1.t6 VB_A.t52 m1m2.t523 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X838 m9m10.t226 bias1.t662 VCC.t498 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X839 VCC.t505 bias1.t663 m1m2.t240 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X840 dummy_9.t185 bias1.t664 dummy_9.t184 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X841 dummy_100.t15 IB.t23 dummy_100.t14 VCC.t7 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X842 dummy_9.t183 bias1.t665 dummy_9.t182 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X843 m9m10.t225 bias1.t666 VCC.t503 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X844 m9m10.t224 bias1.t667 VCC.t504 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X845 VCC.t502 bias1.t668 m1m2.t239 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X846 dummy_9.t181 bias1.t669 dummy_9.t180 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X847 dummy_9.t179 bias1.t670 dummy_9.t178 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X848 m9m10.t223 bias1.t671 VCC.t500 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X849 VCC.t501 bias1.t672 m1m2.t238 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X850 dummy_9.t177 bias1.t57 dummy_9.t176 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X851 VCC.t497 bias1.t673 m1m2.t237 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X852 m9m10.t222 bias1.t674 VCC.t496 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X853 VCC.t495 bias1.t675 m1m2.t236 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X854 dummy_2.t41 VB_A.t53 dummy_2.t40 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X855 m11m12.t13 VB_B.t54 OUT.t57 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X856 VCC.t494 bias1.t676 m1m2.t235 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X857 bias3.t9 IN_M.t19 a_46836_49340.t26 VCC.t9 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X858 m9m10.t221 bias1.t677 VCC.t493 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X859 dummy_9.t175 bias1.t678 dummy_9.t174 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X860 dummy_9.t173 bias1.t679 dummy_9.t172 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X861 VCC.t492 bias1.t680 m1m2.t234 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X862 m9m10.t220 bias1.t681 VCC.t486 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X863 m9m10.t219 bias1.t682 VCC.t485 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X864 VCC.t487 bias1.t683 m1m2.t233 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X865 m9m10.t218 bias1.t684 VCC.t491 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X866 bias21.t3 bias21.t2 VSS.t19 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X867 VCC.t490 bias1.t685 m1m2.t232 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X868 a_46836_49340.t60 IN_P.t16 bias21.t21 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X869 dummy_3.t27 VB_B.t55 dummy_3.t26 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X870 VCC.t489 bias1.t686 m1m2.t231 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X871 dummy_9.t171 bias1.t687 dummy_9.t170 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X872 dummy_2.t39 VB_A.t54 dummy_2.t38 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X873 OUT.t36 VB_B.t56 m11m12.t12 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X874 VCC.t488 bias1.t688 m1m2.t230 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X875 dummy_9.t169 bias1.t57 dummy_9.t168 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X876 VCC.t484 bias1.t689 m1m2.t229 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X877 m9m10.t217 bias1.t690 VCC.t483 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X878 m9m10.t216 bias1.t691 VCC.t482 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X879 m9m10.t215 bias1.t692 VCC.t481 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X880 VCC.t480 bias1.t693 m1m2.t228 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X881 dummy_9.t167 bias1.t694 dummy_9.t166 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X882 VCC.t479 bias1.t695 m1m2.t227 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X883 VCC.t478 bias1.t696 m1m2.t226 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X884 m9m10.t214 bias1.t697 VCC.t476 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X885 VCC.t477 bias1.t698 m1m2.t225 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X886 VCC.t475 bias1.t699 m1m2.t224 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X887 OUT.t15 VB_A.t55 m9m10.t526 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X888 m1m2.t522 VB_A.t56 bias1.t6 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X889 bias1.t0 VB_B.t57 m3m4.t19 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X890 m9m10.t213 bias1.t700 VCC.t474 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X891 VCC.t473 bias1.t701 m1m2.t223 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X892 m9m10.t212 bias1.t702 VCC.t467 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X893 VCC.t472 bias1.t703 m1m2.t222 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X894 dummy_9.t165 bias1.t704 dummy_9.t164 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X895 VCC.t471 bias1.t705 m1m2.t221 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X896 dummy_3.t25 VB_B.t58 dummy_3.t24 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X897 m9m10.t211 bias1.t706 VCC.t470 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X898 VCC.t469 bias1.t707 m1m2.t220 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X899 dummy_9.t163 bias1.t57 dummy_9.t162 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X900 OUT.t14 VB_A.t57 m9m10.t523 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X901 m9m10.t210 bias1.t708 VCC.t468 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X902 m9m10.t209 bias1.t709 VCC.t466 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X903 VCC.t465 bias1.t710 m1m2.t219 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X904 m9m10.t208 bias1.t711 VCC.t464 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X905 dummy_9.t161 bias1.t712 dummy_9.t160 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X906 m9m10.t207 bias1.t713 VCC.t463 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X907 m9m10.t206 bias1.t714 VCC.t462 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X908 VCC.t461 bias1.t715 m1m2.t218 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X909 m9m10.t524 VB_A.t58 OUT.t13 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X910 OUT.t53 VB_B.t59 m11m12.t11 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X911 m9m10.t205 bias1.t716 VCC.t460 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X912 VCC.t459 bias1.t717 m1m2.t217 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X913 VCC.t458 bias1.t718 m1m2.t216 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X914 VCC.t454 bias1.t719 m1m2.t215 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X915 m9m10.t204 bias1.t720 VCC.t457 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X916 VCC.t456 bias1.t721 m1m2.t214 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X917 m3m4.t18 VB_B.t60 bias1.t3 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X918 dummy_9.t159 bias1.t722 dummy_9.t158 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X919 OUT.t12 VB_A.t59 m9m10.t525 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X920 dummy_2.t37 VB_A.t60 dummy_2.t36 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X921 VCC.t455 bias1.t723 m1m2.t213 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X922 dummy_9.t157 bias1.t724 dummy_9.t156 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X923 dummy_9.t155 bias1.t725 dummy_9.t154 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X924 VCC.t453 bias1.t726 m1m2.t212 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X925 m9m10.t203 bias1.t727 VCC.t452 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X926 dummy_9.t153 bias1.t728 dummy_9.t152 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X927 VCC.t451 bias1.t729 m1m2.t211 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X928 VCC.t450 bias1.t730 m1m2.t210 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X929 VCC.t449 bias1.t731 m1m2.t209 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X930 VCC.t447 bias1.t732 m1m2.t208 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X931 m11m12.t10 VB_B.t61 OUT.t33 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X932 dummy_3.t23 VB_B.t62 dummy_3.t22 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X933 VCC.t448 bias1.t733 m1m2.t207 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X934 VCC.t446 bias1.t734 m1m2.t206 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X935 dummy_9.t151 bias1.t735 dummy_9.t150 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X936 m9m10.t202 bias1.t736 VCC.t445 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X937 m9m10.t201 bias1.t737 VCC.t444 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X938 m9m10.t200 bias1.t738 VCC.t443 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X939 VCC.t442 bias1.t739 m1m2.t205 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X940 VCC.t441 bias1.t740 m1m2.t204 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X941 m9m10.t199 bias1.t741 VCC.t440 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X942 m9m10.t198 bias1.t742 VCC.t439 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X943 VCC.t438 bias1.t743 m1m2.t203 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X944 m9m10.t197 bias1.t744 VCC.t437 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X945 VCC.t436 bias1.t745 m1m2.t202 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X946 dummy_9.t149 bias1.t746 dummy_9.t148 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X947 m9m10.t196 bias1.t747 VCC.t435 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X948 m9m10.t195 bias1.t748 VCC.t434 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X949 m9m10.t194 bias1.t749 VCC.t433 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X950 m9m10.t193 bias1.t750 VCC.t432 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X951 m9m10.t192 bias1.t751 VCC.t431 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X952 OUT.t43 VB_B.t63 m11m12.t9 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X953 dummy_9.t147 bias1.t752 dummy_9.t146 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X954 VCC.t430 bias1.t753 m1m2.t201 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X955 VCC.t429 bias1.t754 m1m2.t200 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X956 VCC.t420 bias1.t755 m1m2.t199 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X957 VCC.t428 bias1.t756 m1m2.t198 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X958 m9m10.t191 bias1.t757 VCC.t427 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X959 bias21.t20 IN_P.t17 a_46836_49340.t61 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X960 m9m10.t190 bias1.t758 VCC.t426 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X961 VCC.t421 bias1.t759 m1m2.t197 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X962 bias21.t19 IN_P.t18 a_46836_49340.t14 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X963 m11m12.t30 bias21.t38 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=1
**devattr s=58000,2116 d=58000,2116
X964 VCC.t424 bias1.t760 m1m2.t196 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X965 m9m10.t189 bias1.t761 VCC.t425 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X966 m9m10.t188 bias1.t762 VCC.t423 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X967 dummy_2.t35 VB_A.t61 dummy_2.t34 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X968 dummy_9.t145 bias1.t763 dummy_9.t144 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X969 dummy_9.t143 bias1.t764 dummy_9.t142 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X970 m3m4.t17 VB_B.t64 bias1.t5 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X971 VCC.t422 bias1.t765 m1m2.t195 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X972 VCC.t419 bias1.t766 m1m2.t194 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X973 m9m10.t187 bias1.t767 VCC.t418 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X974 m9m10.t186 bias1.t768 VCC.t417 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X975 dummy_3.t21 VB_B.t65 dummy_3.t20 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X976 bias1.t6 VB_A.t62 m1m2.t520 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X977 VCC.t416 bias1.t769 m1m2.t193 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X978 VCC.t415 bias1.t770 m1m2.t192 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X979 VCC.t414 bias1.t771 m1m2.t191 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X980 VCC.t413 bias1.t772 m1m2.t190 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X981 VCC.t412 bias1.t773 m1m2.t189 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X982 m9m10.t185 bias1.t774 VCC.t411 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X983 m9m10.t184 bias1.t775 VCC.t410 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X984 VCC.t409 bias1.t776 m1m2.t188 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X985 m9m10.t183 bias1.t777 VCC.t408 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X986 m9m10.t182 bias1.t778 VCC.t407 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X987 m9m10.t181 bias1.t779 VCC.t406 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X988 m9m10.t180 bias1.t780 VCC.t404 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X989 m9m10.t179 bias1.t781 VCC.t405 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X990 VCC.t403 bias1.t782 m1m2.t187 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X991 m9m10.t178 bias1.t783 VCC.t402 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X992 VCC.t1048 IB.t2 IB.t3 VCC.t1038 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X993 VCC.t401 bias1.t784 m1m2.t186 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X994 VCC.t400 bias1.t785 m1m2.t185 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X995 VCC.t388 bias1.t786 m1m2.t184 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X996 a_46836_49340.t25 IN_M.t20 bias3.t10 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X997 VCC.t1049 IB.t0 IB.t1 VCC.t1038 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X998 m9m10.t177 bias1.t787 VCC.t399 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X999 bias1.t6 VB_A.t63 m1m2.t517 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1000 dummy_9.t141 bias1.t788 dummy_9.t140 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1001 m9m10.t176 bias1.t789 VCC.t398 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1002 dummy_2.t33 VB_A.t64 dummy_2.t32 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1003 dummy_3.t19 VB_B.t66 dummy_3.t18 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1004 dummy_9.t139 bias1.t790 dummy_9.t138 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1005 m9m10.t175 bias1.t791 VCC.t397 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1006 VCC.t396 bias1.t792 m1m2.t183 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1007 m9m10.t174 bias1.t793 VCC.t395 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1008 VCC.t386 bias1.t794 m1m2.t182 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1009 VCC.t394 bias1.t795 m1m2.t181 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1010 m9m10.t173 bias1.t796 VCC.t393 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1011 VCC.t392 bias1.t797 m1m2.t180 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1012 m9m10.t172 bias1.t798 VCC.t391 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1013 VCC.t387 bias1.t799 m1m2.t179 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1014 VCC.t390 bias1.t800 m1m2.t178 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1015 VCC.t389 bias1.t801 m1m2.t177 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1016 bias21.t18 IN_P.t19 a_46836_49340.t15 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1017 m9m10.t171 bias1.t802 VCC.t385 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1018 dummy_9.t137 bias1.t803 dummy_9.t136 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1019 VCC.t384 bias1.t804 m1m2.t176 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1020 VCC.t382 bias1.t805 m1m2.t175 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1021 m9m10.t170 bias1.t806 VCC.t383 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1022 dummy_9.t135 bias1.t807 dummy_9.t134 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1023 m9m10.t169 bias1.t808 VCC.t381 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1024 VCC.t377 bias1.t809 m1m2.t174 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1025 m9m10.t168 bias1.t810 VCC.t380 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1026 m9m10.t167 bias1.t811 VCC.t379 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1027 VCC.t378 bias1.t812 m1m2.t173 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1028 VCC.t376 bias1.t813 m1m2.t172 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1029 OUT.t50 VB_B.t67 m11m12.t8 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1030 dummy_9.t133 bias1.t814 dummy_9.t132 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1031 VCC.t375 bias1.t815 m1m2.t171 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1032 bias1.t5 VB_B.t68 m3m4.t16 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1033 dummy_3.t17 VB_B.t69 dummy_3.t16 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1034 VCC.t374 bias1.t816 m1m2.t170 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1035 VCC.t373 bias1.t817 m1m2.t169 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1036 m9m10.t166 bias1.t818 VCC.t372 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1037 m9m10.t165 bias1.t819 VCC.t371 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1038 VCC.t370 bias1.t820 m1m2.t168 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1039 m9m10.t164 bias1.t821 VCC.t369 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1040 m9m10.t163 bias1.t822 VCC.t368 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1041 VCC.t367 bias1.t823 m1m2.t167 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1042 m1m2.t518 VB_A.t65 bias1.t6 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1043 VCC.t366 bias1.t824 m1m2.t166 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1044 VCC.t365 bias1.t825 m1m2.t165 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1045 VCC.t364 bias1.t826 m1m2.t164 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1046 m9m10.t162 bias1.t827 VCC.t363 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1047 m9m10.t161 bias1.t828 VCC.t362 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1048 dummy_9.t131 bias1.t829 dummy_9.t130 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1049 OUT.t11 VB_A.t66 m9m10.t519 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1050 dummy_2.t31 VB_A.t67 dummy_2.t30 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1051 m3m4.t15 VB_B.t70 bias1.t5 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1052 m9m10.t160 bias1.t830 VCC.t361 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1053 dummy_100.t13 IB.t24 dummy_100.t12 VCC.t0 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X1054 dummy_3.t15 VB_B.t71 dummy_3.t14 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1055 VCC.t360 bias1.t831 m1m2.t163 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1056 m9m10.t159 bias1.t832 VCC.t359 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1057 VCC.t358 bias1.t833 m1m2.t162 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1058 dummy_9.t129 bias1.t834 dummy_9.t128 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1059 VCC.t357 bias1.t835 m1m2.t161 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1060 VCC.t356 bias1.t836 m1m2.t160 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1061 dummy_4.t19 bias3.t49 dummy_4.t18 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X1062 m9m10.t158 bias1.t837 VCC.t16 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1063 VCC.t355 bias1.t838 m1m2.t159 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1064 dummy_9.t127 bias1.t231 dummy_9.t126 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1065 m9m10.t157 bias1.t839 VCC.t18 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1066 VCC.t354 bias1.t840 m1m2.t158 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1067 VCC.t33 bias1.t841 m1m2.t157 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1068 m9m10.t156 bias1.t842 VCC.t353 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1069 dummy_100.t11 IB.t25 dummy_100.t10 VCC.t1038 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X1070 dummy_100.t9 IB.t26 dummy_100.t8 VCC.t6 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X1071 m9m10.t155 bias1.t843 VCC.t352 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1072 VCC.t351 bias1.t844 m1m2.t156 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1073 dummy_9.t125 bias1.t845 dummy_9.t124 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1074 VCC.t350 bias1.t846 m1m2.t155 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1075 VCC.t349 bias1.t847 m1m2.t154 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1076 m9m10.t154 bias1.t848 VCC.t348 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1077 dummy_4.t17 bias3.t50 dummy_4.t16 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X1078 m9m10.t153 bias1.t849 VCC.t347 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1079 dummy_9.t123 bias1.t850 dummy_9.t122 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1080 m1m2.t514 VB_A.t68 bias1.t6 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1081 VCC.t346 bias1.t851 m1m2.t153 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1082 VCC.t345 bias1.t852 m1m2.t152 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1083 VCC.t344 bias1.t853 m1m2.t151 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1084 dummy_2.t29 VB_A.t69 dummy_2.t28 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1085 bias1.t2 VB_B.t72 m3m4.t14 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1086 m9m10.t152 bias1.t854 VCC.t343 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1087 VCC.t342 bias1.t855 m1m2.t150 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1088 VCC.t341 bias1.t856 m1m2.t149 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1089 m9m10.t151 bias1.t857 VCC.t340 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1090 VCC.t339 bias1.t858 m1m2.t148 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1091 dummy_9.t121 bias1.t859 dummy_9.t120 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1092 dummy_2.t27 VB_A.t70 dummy_2.t26 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1093 dummy_2.t25 VB_A.t71 dummy_2.t24 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1094 dummy_3.t13 VB_B.t73 dummy_3.t12 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1095 dummy_9.t119 bias1.t860 dummy_9.t118 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1096 dummy_9.t117 bias1.t861 dummy_9.t116 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1097 bias1.t4 VB_B.t74 m3m4.t13 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1098 VCC.t338 bias1.t862 m1m2.t147 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1099 m9m10.t150 bias1.t863 VCC.t337 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1100 VCC.t336 bias1.t864 m1m2.t146 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1101 m9m10.t149 bias1.t865 VCC.t335 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1102 VCC.t334 bias1.t866 m1m2.t145 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1103 dummy_9.t115 bias1.t867 dummy_9.t114 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1104 VCC.t333 bias1.t868 m1m2.t144 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1105 VCC.t332 bias1.t869 m1m2.t143 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1106 m9m10.t148 bias1.t870 VCC.t331 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1107 m1m2.t512 VB_A.t72 bias1.t6 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1108 dummy_2.t23 VB_A.t73 dummy_2.t22 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1109 m9m10.t147 bias1.t871 VCC.t330 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1110 m9m10.t146 bias1.t872 VCC.t329 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1111 dummy_9.t113 bias1.t873 dummy_9.t112 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1112 VCC.t325 bias1.t874 m1m2.t142 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1113 VCC.t328 bias1.t875 m1m2.t141 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1114 VCC.t327 bias1.t876 m1m2.t140 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1115 VCC.t326 bias1.t877 m1m2.t139 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1116 m9m10.t145 bias1.t878 VCC.t324 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1117 VCC.t323 bias1.t879 m1m2.t138 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1118 dummy_9.t111 bias1.t880 dummy_9.t110 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1119 VCC.t322 bias1.t881 m1m2.t137 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1120 a_46836_49340.t24 IN_M.t21 bias3.t11 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1121 dummy_4.t15 bias3.t51 dummy_4.t14 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X1122 m9m10.t144 bias1.t882 VCC.t321 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1123 VCC.t320 bias1.t883 m1m2.t136 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1124 m9m10.t143 bias1.t884 VCC.t319 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1125 m9m10.t142 bias1.t885 VCC.t318 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1126 VCC.t317 bias1.t886 m1m2.t135 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1127 dummy_9.t109 bias1.t887 dummy_9.t108 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1128 bias3.t24 IN_M.t22 a_46836_49340.t23 VCC.t9 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1129 dummy_100.t7 IB.t27 dummy_100.t6 VCC.t6 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X1130 m9m10.t141 bias1.t888 VCC.t316 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1131 m9m10.t140 bias1.t889 VCC.t315 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1132 VCC.t314 bias1.t890 m1m2.t134 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1133 dummy_9.t107 bias1.t891 dummy_9.t106 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1134 bias1.t1 VB_B.t75 m3m4.t12 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1135 VSS.t15 bias3.t0 bias3.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X1136 m9m10.t139 bias1.t892 VCC.t313 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1137 dummy_9.t105 bias1.t893 dummy_9.t104 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1138 m9m10.t138 bias1.t894 VCC.t312 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1139 VCC.t311 bias1.t895 m1m2.t133 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1140 bias1.t1 VB_B.t76 m3m4.t11 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1141 VCC.t310 bias1.t896 m1m2.t132 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1142 m9m10.t516 VB_A.t74 OUT.t10 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1143 m9m10.t137 bias1.t897 VCC.t309 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1144 dummy_9.t103 bias1.t898 dummy_9.t102 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1145 m9m10.t136 bias1.t899 VCC.t308 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1146 dummy_100.t5 IB.t28 dummy_100.t4 VCC.t8 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X1147 m9m10.t135 bias1.t900 VCC.t307 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1148 VCC.t306 bias1.t901 m1m2.t131 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1149 VCC.t305 bias1.t902 m1m2.t130 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1150 dummy_9.t101 bias1.t903 dummy_9.t100 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1151 dummy_9.t99 bias1.t904 dummy_9.t98 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1152 dummy_9.t97 bias1.t905 dummy_9.t96 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1153 dummy_9.t95 bias1.t906 dummy_9.t94 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1154 VCC.t304 bias1.t907 m1m2.t129 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1155 m9m10.t134 bias1.t908 VCC.t303 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1156 VCC.t23 bias1.t909 m1m2.t128 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1157 m9m10.t133 bias1.t910 VCC.t302 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1158 VCC.t301 bias1.t911 m1m2.t127 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1159 VCC.t300 bias1.t912 m1m2.t126 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1160 m9m10.t132 bias1.t913 VCC.t299 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1161 VCC.t298 bias1.t914 m1m2.t125 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1162 VCC.t27 bias1.t915 m1m2.t124 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1163 m9m10.t131 bias1.t916 VCC.t36 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1164 VCC.t297 bias1.t917 m1m2.t123 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1165 VCC.t38 bias1.t918 m1m2.t122 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1166 m9m10.t130 bias1.t919 VCC.t296 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1167 m9m10.t129 bias1.t920 VCC.t295 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1168 dummy_9.t93 bias1.t921 dummy_9.t92 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1169 VCC.t294 bias1.t922 m1m2.t121 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1170 a_46836_49340.t64 IN_P.t20 bias21.t17 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1171 m9m10.t128 bias1.t923 VCC.t267 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1172 VCC.t293 bias1.t924 m1m2.t120 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1173 m9m10.t127 bias1.t925 VCC.t292 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1174 VCC.t291 bias1.t926 m1m2.t119 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1175 a_46836_49340.t22 IN_M.t23 bias3.t25 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1176 dummy_4.t13 bias3.t52 dummy_4.t12 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X1177 VCC.t290 bias1.t927 m1m2.t118 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1178 VCC.t289 bias1.t928 m1m2.t117 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1179 m9m10.t126 bias1.t929 VCC.t288 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1180 bias1.t4 VB_B.t77 m3m4.t10 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1181 dummy_9.t91 bias1.t930 dummy_9.t90 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1182 dummy_2.t21 VB_A.t75 dummy_2.t20 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1183 m9m10.t125 bias1.t931 VCC.t287 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1184 VCC.t266 bias1.t932 m1m2.t116 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1185 dummy_9.t89 bias1.t933 dummy_9.t88 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1186 m9m10.t124 bias1.t934 VCC.t286 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1187 VCC.t285 bias1.t935 m1m2.t115 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1188 m9m10.t123 bias1.t936 VCC.t284 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1189 VCC.t268 bias1.t937 m1m2.t114 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1190 m9m10.t122 bias1.t938 VCC.t283 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1191 m9m10.t121 bias1.t939 VCC.t282 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1192 a_46836_49340.t65 IN_P.t21 bias21.t16 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1193 VCC.t281 bias1.t940 m1m2.t113 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1194 m9m10.t120 bias1.t941 VCC.t280 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1195 OUT.t47 VB_B.t78 m11m12.t7 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1196 dummy_9.t87 bias1.t942 dummy_9.t86 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1197 m9m10.t119 bias1.t943 VCC.t279 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1198 VCC.t278 bias1.t944 m1m2.t112 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1199 VCC.t277 bias1.t945 m1m2.t111 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1200 m9m10.t118 bias1.t946 VCC.t276 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1201 VCC.t275 bias1.t947 m1m2.t110 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1202 bias1.t1 VB_B.t79 m3m4.t9 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1203 dummy_4.t11 bias3.t53 dummy_4.t10 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X1204 VCC.t272 bias1.t948 m1m2.t109 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1205 VCC.t273 bias1.t949 m1m2.t108 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1206 m9m10.t117 bias1.t950 VCC.t274 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1207 m3m4.t8 VB_B.t80 bias1.t5 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1208 VCC.t271 bias1.t951 m1m2.t107 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1209 m9m10.t116 bias1.t952 VCC.t270 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1210 m9m10.t115 bias1.t953 VCC.t269 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1211 VCC.t265 bias1.t954 m1m2.t106 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1212 dummy_9.t85 bias1.t955 dummy_9.t84 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1213 VCC.t264 bias1.t956 m1m2.t105 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1214 m9m10.t114 bias1.t957 VCC.t263 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1215 a_46836_49340.t4 IN_P.t22 bias21.t15 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1216 m9m10.t113 bias1.t958 VCC.t262 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1217 VCC.t261 bias1.t959 m1m2.t104 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1218 OUT.t9 VB_A.t76 m9m10.t513 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1219 m1m2.t511 VB_A.t77 bias1.t6 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1220 VCC.t257 bias1.t960 m1m2.t103 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1221 m9m10.t112 bias1.t961 VCC.t260 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1222 m9m10.t111 bias1.t962 VCC.t259 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1223 VCC.t258 bias1.t963 m1m2.t102 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1224 m9m10.t110 bias1.t964 VCC.t256 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1225 VCC.t255 bias1.t965 m1m2.t101 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1226 VCC.t254 bias1.t966 m1m2.t100 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1227 m9m10.t109 bias1.t967 VCC.t253 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1228 a_46836_49340.t48 IB.t29 VCC.t1037 VCC.t0 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X1229 m9m10.t108 bias1.t968 VCC.t252 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1230 a_46836_49340.t47 IB.t30 VCC.t1045 VCC.t0 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X1231 VCC.t177 bias1.t969 m1m2.t99 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1232 VCC.t251 bias1.t970 m1m2.t98 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1233 m9m10.t107 bias1.t971 VCC.t250 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1234 m9m10.t106 bias1.t972 VCC.t178 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1235 m9m10.t105 bias1.t973 VCC.t249 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1236 dummy_9.t83 bias1.t974 dummy_9.t82 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1237 VCC.t248 bias1.t975 m1m2.t97 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1238 VCC.t247 bias1.t976 m1m2.t96 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1239 VCC.t246 bias1.t977 m1m2.t95 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1240 VCC.t245 bias1.t978 m1m2.t94 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1241 m9m10.t104 bias1.t979 VCC.t244 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1242 bias1.t6 VB_A.t78 m1m2.t508 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1243 m3m4.t7 VB_B.t81 bias1.t2 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1244 m9m10.t103 bias1.t980 VCC.t243 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1245 OUT.t8 VB_A.t79 m9m10.t512 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1246 VCC.t242 bias1.t981 m1m2.t93 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1247 dummy_2.t19 VB_A.t80 dummy_2.t18 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1248 VCC.t240 bias1.t982 m1m2.t92 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1249 m9m10.t102 bias1.t983 VCC.t241 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1250 bias1.t3 VB_B.t82 m3m4.t6 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1251 VCC.t239 bias1.t984 m1m2.t91 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1252 dummy_9.t81 bias1.t985 dummy_9.t80 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1253 dummy_2.t17 VB_A.t81 dummy_2.t16 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1254 m9m10.t101 bias1.t986 VCC.t238 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1255 m11m12.t6 VB_B.t83 OUT.t34 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1256 VCC.t175 bias1.t987 m1m2.t90 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1257 m9m10.t100 bias1.t988 VCC.t237 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1258 m9m10.t99 bias1.t989 VCC.t236 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1259 m9m10.t98 bias1.t990 VCC.t179 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1260 VCC.t235 bias1.t991 m1m2.t89 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1261 dummy_9.t79 bias1.t992 dummy_9.t78 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1262 VCC.t234 bias1.t993 m1m2.t88 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1263 m9m10.t97 bias1.t994 VCC.t233 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1264 dummy_3.t11 VB_B.t84 dummy_3.t10 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1265 OUT.t7 VB_A.t82 m9m10.t510 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1266 m1m2.t507 VB_A.t83 bias1.t6 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1267 dummy_2.t15 VB_A.t84 dummy_2.t14 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1268 m9m10.t96 bias1.t995 VCC.t232 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1269 VCC.t231 bias1.t996 m1m2.t87 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1270 m9m10.t95 bias1.t997 VCC.t230 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1271 OUT.t35 VB_B.t85 m11m12.t5 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1272 dummy_9.t77 bias1.t998 dummy_9.t76 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1273 m9m10.t94 bias1.t999 VCC.t222 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1274 VCC.t229 bias1.t1000 m1m2.t86 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1275 m9m10.t93 bias1.t1001 VCC.t228 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1276 m9m10.t92 bias1.t1002 VCC.t227 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1277 dummy_4.t9 bias3.t54 dummy_4.t8 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X1278 dummy_9.t75 bias1.t1003 dummy_9.t74 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1279 VCC.t226 bias1.t1004 m1m2.t85 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1280 m9m10.t91 bias1.t1005 VCC.t225 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1281 VCC.t224 bias1.t1006 m1m2.t84 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1282 a_46836_49340.t5 IN_P.t23 bias21.t14 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1283 m9m10.t90 bias1.t1007 VCC.t223 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1284 VCC.t221 bias1.t1008 m1m2.t83 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1285 dummy_9.t73 bias1.t231 dummy_9.t72 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1286 VCC.t220 bias1.t1009 m1m2.t82 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1287 m9m10.t89 bias1.t1010 VCC.t219 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1288 bias21.t13 IN_P.t24 a_46836_49340.t52 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1289 m9m10.t507 VB_A.t85 OUT.t6 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1290 m9m10.t88 bias1.t1011 VCC.t218 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1291 VCC.t207 bias1.t1012 m1m2.t81 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1292 m9m10.t87 bias1.t1013 VCC.t217 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1293 dummy_9.t71 bias1.t1014 dummy_9.t70 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1294 m9m10.t86 bias1.t1015 VCC.t208 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1295 m9m10.t85 bias1.t1016 VCC.t216 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1296 m3m4.t5 VB_B.t86 bias1.t1 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1297 VCC.t209 bias1.t1017 m1m2.t80 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1298 dummy_9.t69 bias1.t1018 dummy_9.t68 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1299 VCC.t1046 IB.t31 a_46836_49340.t46 VCC.t2 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X1300 m9m10.t84 bias1.t1019 VCC.t215 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1301 VCC.t214 bias1.t1020 m1m2.t79 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1302 VCC.t213 bias1.t1021 m1m2.t78 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1303 m11m12.t4 VB_B.t87 OUT.t46 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1304 m9m10.t83 bias1.t1022 VCC.t212 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1305 VCC.t211 bias1.t1023 m1m2.t77 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1306 m9m10.t508 VB_A.t86 OUT.t5 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1307 m9m10.t82 bias1.t1024 VCC.t210 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1308 m9m10.t81 bias1.t1025 VCC.t206 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1309 m9m10.t80 bias1.t1026 VCC.t205 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1310 VCC.t204 bias1.t1027 m1m2.t76 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1311 m9m10.t79 bias1.t1028 VCC.t203 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1312 dummy_9.t67 bias1.t1029 dummy_9.t66 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1313 VCC.t202 bias1.t1030 m1m2.t75 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1314 dummy_9.t65 bias1.t1031 dummy_9.t64 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1315 dummy_9.t63 bias1.t1032 dummy_9.t62 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1316 VCC.t201 bias1.t1033 m1m2.t74 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1317 m9m10.t78 bias1.t1034 VCC.t200 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1318 m9m10.t77 bias1.t1035 VCC.t199 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1319 dummy_9.t61 bias1.t1036 dummy_9.t60 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1320 m9m10.t76 bias1.t1037 VCC.t198 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1321 VCC.t197 bias1.t1038 m1m2.t73 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1322 m9m10.t75 bias1.t1039 VCC.t196 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1323 m9m10.t505 VB_A.t87 OUT.t4 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1324 m9m10.t74 bias1.t1040 VCC.t195 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1325 dummy_9.t59 bias1.t1041 dummy_9.t58 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1326 m9m10.t73 bias1.t1042 VCC.t21 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1327 dummy_9.t57 bias1.t1043 dummy_9.t56 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1328 VCC.t194 bias1.t1044 m1m2.t72 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1329 m9m10.t72 bias1.t1045 VCC.t19 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1330 VCC.t176 bias1.t1046 m1m2.t71 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1331 VCC.t193 bias1.t1047 m1m2.t70 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1332 m9m10.t71 bias1.t1048 VCC.t192 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1333 VCC.t191 bias1.t1049 m1m2.t69 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1334 bias1.t3 VB_B.t88 m3m4.t4 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1335 VCC.t190 bias1.t1050 m1m2.t68 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1336 a_46836_49340.t53 IN_P.t25 bias21.t12 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1337 m9m10.t70 bias1.t1051 VCC.t189 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1338 VCC.t188 bias1.t1052 m1m2.t67 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1339 m9m10.t69 bias1.t1053 VCC.t187 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1340 dummy_2.t13 VB_A.t88 dummy_2.t12 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1341 bias3.t22 IN_M.t24 a_46836_49340.t21 VCC.t9 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1342 m9m10.t68 bias1.t1054 VCC.t186 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1343 dummy_9.t55 bias1.t1055 dummy_9.t54 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1344 m11m12.t3 VB_B.t89 OUT.t45 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1345 m9m10.t67 bias1.t1056 VCC.t185 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1346 VCC.t184 bias1.t1057 m1m2.t66 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1347 dummy_2.t11 VB_A.t89 dummy_2.t10 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1348 dummy_9.t53 bias1.t1058 dummy_9.t52 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1349 VCC.t183 bias1.t1059 m1m2.t65 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1350 dummy_9.t51 bias1.t1060 dummy_9.t50 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1351 m9m10.t66 bias1.t1061 VCC.t182 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1352 VCC.t181 bias1.t1062 m1m2.t64 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1353 m9m10.t65 bias1.t1063 VCC.t180 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1354 m9m10.t64 bias1.t1064 VCC.t174 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1355 VCC.t25 bias1.t1065 m1m2.t63 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1356 dummy_9.t49 bias1.t1066 dummy_9.t48 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1357 m9m10.t63 bias1.t1067 VCC.t173 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1358 m1m2.t503 VB_A.t90 bias1.t6 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1359 VCC.t172 bias1.t1068 m1m2.t62 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1360 dummy_3.t9 VB_B.t90 dummy_3.t8 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1361 VCC.t168 bias1.t1069 m1m2.t61 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1362 m9m10.t62 bias1.t1070 VCC.t170 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1363 VCC.t171 bias1.t1071 m1m2.t60 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1364 dummy_9.t47 bias1.t1072 dummy_9.t46 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1365 bias1.t2 VB_B.t91 m3m4.t3 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1366 m9m10.t61 bias1.t1073 VCC.t169 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1367 VCC.t167 bias1.t1074 m1m2.t59 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1368 dummy_9.t45 bias1.t1075 dummy_9.t44 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1369 VCC.t166 bias1.t1076 m1m2.t58 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1370 m9m10.t60 bias1.t1077 VCC.t165 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1371 dummy_4.t7 bias3.t55 dummy_4.t6 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X1372 VCC.t164 bias1.t1078 m1m2.t57 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1373 m9m10.t59 bias1.t1079 VCC.t163 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1374 VCC.t162 bias1.t1080 m1m2.t56 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1375 m9m10.t58 bias1.t1081 VCC.t161 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1376 VCC.t160 bias1.t1082 m1m2.t55 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1377 m9m10.t57 bias1.t1083 VCC.t159 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1378 dummy_9.t43 bias1.t1084 dummy_9.t42 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1379 m3m4.t2 VB_B.t92 bias1.t1 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1380 VCC.t158 bias1.t1085 m1m2.t54 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1381 dummy_4.t5 bias3.t56 dummy_4.t4 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X1382 m9m10.t56 bias1.t1086 VCC.t157 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1383 VCC.t155 bias1.t1087 m1m2.t53 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1384 m9m10.t55 bias1.t1088 VCC.t156 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1385 m9m10.t54 bias1.t1089 VCC.t154 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1386 VCC.t153 bias1.t1090 m1m2.t52 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1387 VCC.t152 bias1.t1091 m1m2.t51 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1388 VCC.t151 bias1.t1092 m1m2.t50 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1389 dummy_3.t7 VB_B.t93 dummy_3.t6 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1390 VCC.t147 bias1.t1093 m1m2.t49 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1391 m9m10.t53 bias1.t1094 VCC.t150 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1392 m9m10.t52 bias1.t1095 VCC.t149 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1393 dummy_9.t41 bias1.t1096 dummy_9.t40 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1394 m9m10.t51 bias1.t1097 VCC.t148 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1395 m9m10.t50 bias1.t1098 VCC.t146 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1396 VCC.t145 bias1.t1099 m1m2.t48 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1397 OUT.t3 VB_A.t91 m9m10.t503 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1398 VCC.t143 bias1.t1100 m1m2.t47 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1399 m9m10.t49 bias1.t1101 VCC.t144 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1400 m9m10.t48 bias1.t1102 VCC.t142 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1401 dummy_3.t5 VB_B.t94 dummy_3.t4 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1402 dummy_9.t39 bias1.t1103 dummy_9.t38 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1403 VCC.t141 bias1.t1104 m1m2.t46 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1404 VCC.t110 bias1.t1105 m1m2.t45 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1405 VCC.t140 bias1.t1106 m1m2.t44 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1406 m9m10.t47 bias1.t1107 VCC.t139 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1407 dummy_9.t37 bias1.t207 dummy_9.t36 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1408 dummy_100.t3 IB.t32 dummy_100.t2 VCC.t6 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X1409 m1m2.t504 VB_A.t92 bias1.t6 VCC.t1044 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1410 VCC.t138 bias1.t1108 m1m2.t43 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1411 m9m10.t46 bias1.t1109 VCC.t137 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1412 m11m12.t2 VB_B.t95 OUT.t42 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1413 m9m10.t45 bias1.t1110 VCC.t136 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1414 dummy_2.t9 VB_A.t93 dummy_2.t8 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1415 dummy_9.t35 bias1.t1111 dummy_9.t34 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1416 dummy_9.t33 bias1.t1112 dummy_9.t32 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1417 VCC.t135 bias1.t1113 m1m2.t42 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1418 m9m10.t44 bias1.t1114 VCC.t134 VCC.t133 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1419 m9m10.t43 bias1.t1115 VCC.t132 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1420 dummy_9.t31 bias1.t1116 dummy_9.t30 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1421 m9m10.t42 bias1.t1117 VCC.t131 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1422 dummy_4.t3 bias3.t57 dummy_4.t2 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X1423 VCC.t130 bias1.t1118 m1m2.t41 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1424 VCC.t112 bias1.t1119 m1m2.t40 VCC.t109 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1425 m9m10.t41 bias1.t1120 VCC.t129 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1426 VCC.t128 bias1.t1121 m1m2.t39 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1427 dummy_9.t29 bias1.t1122 dummy_9.t28 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1428 m9m10.t40 bias1.t1123 VCC.t111 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1429 VCC.t113 bias1.t1124 m1m2.t38 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1430 m9m10.t39 bias1.t1125 VCC.t127 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1431 m9m10.t38 bias1.t1126 VCC.t126 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1432 VCC.t125 bias1.t1127 m1m2.t37 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1433 m9m10.t37 bias1.t1128 VCC.t124 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1434 m11m12.t1 VB_B.t96 OUT.t37 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1435 m9m10.t36 bias1.t1129 VCC.t122 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1436 m9m10.t35 bias1.t1130 VCC.t123 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1437 dummy_100.t1 IB.t33 dummy_100.t0 VCC.t6 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=3
**devattr d=58000,2116
X1438 dummy_9.t27 bias1.t1131 dummy_9.t26 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1439 bias21.t1 bias21.t0 VSS.t20 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X1440 VCC.t121 bias1.t1132 m1m2.t36 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1441 m9m10.t34 bias1.t1133 VCC.t120 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1442 VCC.t119 bias1.t1134 m1m2.t35 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1443 dummy_3.t3 VB_B.t97 dummy_3.t2 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1444 m9m10.t33 bias1.t1135 VCC.t118 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1445 m9m10.t32 bias1.t1136 VCC.t116 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1446 VCC.t117 bias1.t1137 m1m2.t34 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1447 VCC.t115 bias1.t1138 m1m2.t33 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1448 m9m10.t31 bias1.t1139 VCC.t114 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1449 m9m10.t30 bias1.t1140 VCC.t108 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1450 VCC.t107 bias1.t1141 m1m2.t32 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1451 OUT.t2 VB_A.t94 m9m10.t502 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1452 bias1.t2 VB_B.t98 m3m4.t1 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1453 m9m10.t29 bias1.t1142 VCC.t106 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1454 VCC.t105 bias1.t1143 m1m2.t31 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1455 dummy_9.t25 bias1.t1144 dummy_9.t24 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1456 m9m10.t28 bias1.t1145 VCC.t104 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1457 VCC.t103 bias1.t1146 m1m2.t30 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1458 VCC.t102 bias1.t1147 m1m2.t29 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1459 m9m10.t27 bias1.t1148 VCC.t98 VCC.t97 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1460 m9m10.t26 bias1.t1149 VCC.t101 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1461 VCC.t100 bias1.t1150 m1m2.t28 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1462 VCC.t99 bias1.t1151 m1m2.t27 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1463 VCC.t96 bias1.t1152 m1m2.t26 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1464 VCC.t95 bias1.t1153 m1m2.t25 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1465 m9m10.t25 bias1.t1154 VCC.t92 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1466 VCC.t93 bias1.t1155 m1m2.t24 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1467 dummy_9.t23 bias1.t207 dummy_9.t22 VCC.t94 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1468 VCC.t91 bias1.t1156 m1m2.t23 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1469 m9m10.t24 bias1.t1157 VCC.t90 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1470 dummy_2.t7 VB_A.t95 dummy_2.t6 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1471 VCC.t89 bias1.t1158 m1m2.t22 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1472 m9m10.t23 bias1.t1159 VCC.t88 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1473 m9m10.t501 VB_A.t96 OUT.t1 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1474 m9m10.t22 bias1.t1160 VCC.t87 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1475 bias3.t23 IN_M.t25 a_46836_49340.t20 VCC.t9 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1476 m9m10.t21 bias1.t1161 VCC.t86 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1477 dummy_9.t21 bias1.t1162 dummy_9.t20 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1478 m9m10.t20 bias1.t1163 VCC.t84 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1479 m9m10.t19 bias1.t1164 VCC.t85 VCC.t17 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1480 VCC.t83 bias1.t1165 m1m2.t21 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1481 dummy_9.t19 bias1.t1166 dummy_9.t18 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1482 VCC.t82 bias1.t1167 m1m2.t20 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1483 a_46836_49340.t8 IN_P.t26 bias21.t11 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1484 m9m10.t18 bias1.t1168 VCC.t81 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1485 bias1.t6 VB_A.t97 m1m2.t500 VCC.t1042 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1486 m9m10.t17 bias1.t1169 VCC.t80 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1487 VCC.t79 bias1.t1170 m1m2.t19 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1488 a_46836_49340.t9 IN_P.t27 bias21.t10 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1489 a_46836_49340.t19 IN_M.t26 bias3.t30 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1490 m9m10.t16 bias1.t1171 VCC.t78 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1491 VCC.t77 bias1.t1172 m1m2.t18 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1492 m9m10.t15 bias1.t1173 VCC.t76 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1493 m9m10.t14 bias1.t1174 VCC.t75 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1494 VCC.t74 bias1.t1175 m1m2.t17 VCC.t73 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1495 dummy_9.t17 bias1.t1176 dummy_9.t16 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1496 dummy_3.t1 VB_B.t99 dummy_3.t0 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1497 VCC.t72 bias1.t1177 m1m2.t16 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1498 VCC.t71 bias1.t1178 m1m2.t15 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1499 m9m10.t13 bias1.t1179 VCC.t70 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1500 VCC.t69 bias1.t1180 m1m2.t14 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1501 VCC.t68 bias1.t1181 m1m2.t13 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1502 m9m10.t12 bias1.t1182 VCC.t67 VCC.t66 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1503 VCC.t65 bias1.t1183 m1m2.t12 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1504 VCC.t64 bias1.t1184 m1m2.t11 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1505 m9m10.t11 bias1.t1185 VCC.t62 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1506 VCC.t63 bias1.t1186 m1m2.t10 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1507 VCC.t61 bias1.t1187 m1m2.t9 VCC.t60 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1508 a_46836_49340.t12 IN_P.t28 bias21.t9 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1509 a_46836_49340.t18 IN_M.t27 bias3.t31 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1510 bias1.t3 VB_B.t100 m3m4.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1511 dummy_2.t5 VB_A.t98 dummy_2.t4 VCC.t1043 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1512 dummy_2.t3 VB_A.t99 dummy_2.t2 VCC.t1039 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1513 VCC.t59 bias1.t1188 m1m2.t8 VCC.t58 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1514 VCC.t57 bias1.t1189 m1m2.t7 VCC.t32 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1515 m9m10.t10 bias1.t1190 VCC.t56 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1516 dummy_9.t15 bias1.t1191 dummy_9.t14 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1517 dummy_9.t13 bias1.t1192 dummy_9.t12 VCC.t55 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1518 dummy_4.t1 bias3.t58 dummy_4.t0 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.25 l=1
**devattr d=14500,616
X1519 m9m10.t9 bias1.t1193 VCC.t54 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1520 dummy_9.t11 bias1.t1194 dummy_9.t10 VCC.t26 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1521 m9m10.t8 bias1.t1195 VCC.t24 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1522 dummy_9.t9 bias1.t1196 dummy_9.t8 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1523 dummy_9.t7 bias1.t1197 dummy_9.t6 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1524 m9m10.t7 bias1.t1198 VCC.t31 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1525 VCC.t53 bias1.t1199 m1m2.t6 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1526 m9m10.t6 bias1.t1200 VCC.t52 VCC.t51 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1527 dummy_9.t5 bias1.t1201 dummy_9.t4 VCC.t37 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1528 VCC.t50 bias1.t1202 m1m2.t5 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1529 bias21.t8 IN_P.t29 a_46836_49340.t13 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1530 m11m12.t0 VB_B.t101 OUT.t38 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1531 VCC.t49 bias1.t1203 m1m2.t4 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1532 m9m10.t5 bias1.t1204 VCC.t48 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1533 dummy_2.t1 VB_A.t100 dummy_2.t0 VCC.t1040 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr d=58000,2116
X1534 bias3.t26 IN_M.t28 a_46836_49340.t17 VCC.t9 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1535 dummy_9.t3 bias1.t1205 dummy_9.t2 VCC.t47 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1536 m9m10.t4 bias1.t1206 VCC.t46 VCC.t45 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1537 dummy_9.t1 bias1.t1207 dummy_9.t0 VCC.t44 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr d=58000,2116
X1538 VCC.t43 bias1.t1208 m1m2.t3 VCC.t42 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1539 VCC.t41 bias1.t1209 m1m2.t2 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1540 m9m10.t3 bias1.t1210 VCC.t30 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1541 m9m10.t2 bias1.t1211 VCC.t29 VCC.t28 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1542 VCC.t35 bias1.t1212 m1m2.t1 VCC.t34 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1543 m9m10.t1 bias1.t1213 VCC.t40 VCC.t15 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1544 VCC.t39 bias1.t1214 m1m2.t0 VCC.t22 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1545 a_46836_49340.t16 IN_M.t29 bias3.t27 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1546 OUT.t0 VB_A.t101 m9m10.t500 VCC.t1041 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1547 m9m10.t0 bias1.t1215 VCC.t14 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=15
**devattr s=58000,2116 d=58000,2116
R0 bias1 bias1.t6 19.8568
R1 bias1.n10 bias1.t829 4.91497
R2 bias1.n10 bias1.t267 4.7605
R3 bias1.n10 bias1.t1162 4.7605
R4 bias1.n10 bias1.t249 4.7605
R5 bias1.n10 bias1.t605 4.7605
R6 bias1.n10 bias1.t378 4.7605
R7 bias1.n10 bias1.t643 4.7605
R8 bias1.n10 bias1.t359 4.7605
R9 bias1.n11 bias1.t903 4.7605
R10 bias1.n11 bias1.t401 4.7605
R11 bias1.n11 bias1.t102 4.7605
R12 bias1.n11 bias1.t665 4.7605
R13 bias1.n11 bias1.t725 4.7605
R14 bias1.n11 bias1.t80 4.7605
R15 bias1.n11 bias1.t763 4.7605
R16 bias1.n11 bias1.t507 4.7605
R17 bias1.n12 bias1.t1029 4.7605
R18 bias1.n12 bias1.t491 4.7605
R19 bias1.n12 bias1.t1072 4.7605
R20 bias1.n12 bias1.t790 4.7605
R21 bias1.n12 bias1.t860 4.7605
R22 bias1.n12 bias1.t233 4.7605
R23 bias1.n12 bias1.t1196 4.7605
R24 bias1.n12 bias1.t281 4.7605
R25 bias1.n13 bias1.t1176 4.7605
R26 bias1.n13 bias1.t620 4.7605
R27 bias1.n13 bias1.t11 4.7605
R28 bias1.n13 bias1.t933 4.7605
R29 bias1.n13 bias1.t654 4.7605
R30 bias1.n13 bias1.t372 4.7605
R31 bias1.n13 bias1.t69 4.7605
R32 bias1.n13 bias1.t417 4.7605
R33 bias1.n14 bias1.t115 4.7605
R34 bias1.n14 bias1.t678 4.7605
R35 bias1.n14 bias1.t100 4.7605
R36 bias1.n14 bias1.t1060 4.7605
R37 bias1.n14 bias1.t1058 4.7605
R38 bias1.n14 bias1.t518 4.7605
R39 bias1.n14 bias1.t1041 4.7605
R40 bias1.n14 bias1.t555 4.7605
R41 bias1.n15 bias1.t269 4.7605
R42 bias1.n15 bias1.t803 4.7605
R43 bias1.n15 bias1.t254 4.7605
R44 bias1.n15 bias1.t845 4.7605
R45 bias1.n15 bias1.t1207 4.7605
R46 bias1.n15 bias1.t645 4.7605
R47 bias1.n15 bias1.t1191 4.7605
R48 bias1.n15 bias1.t905 4.7605
R49 bias1.n16 bias1.t22 4.7605
R50 bias1.n16 bias1.t942 4.7605
R51 bias1.n16 bias1.t388 4.7605
R52 bias1.n16 bias1.t930 4.7605
R53 bias1.n16 bias1.t144 4.7605
R54 bias1.n16 bias1.t426 4.7605
R55 bias1.n16 bias1.t128 4.7605
R56 bias1.n16 bias1.t1032 4.7605
R57 bias1.n17 bias1.t169 4.7605
R58 bias1.n17 bias1.t1075 4.7605
R59 bias1.n17 bias1.t461 4.7605
R60 bias1.n17 bias1.t1055 4.7605
R61 bias1.n17 bias1.t296 4.7605
R62 bias1.n17 bias1.t834 4.7605
R63 bias1.n17 bias1.t283 4.7605
R64 bias1.n17 bias1.t814 4.7605
R65 bias1.n18 bias1.t321 4.7605
R66 bias1.n18 bias1.t14 4.7605
R67 bias1.n18 bias1.t593 4.7605
R68 bias1.n18 bias1.t1205 4.7605
R69 bias1.n18 bias1.t579 4.7605
R70 bias1.n18 bias1.t313 4.7605
R71 bias1.n18 bias1.t921 4.7605
R72 bias1.n18 bias1.t293 4.7605
R73 bias1.n19 bias1.t1197 4.7605
R74 bias1.n19 bias1.t338 4.7605
R75 bias1.n19 bias1.t26 4.7605
R76 bias1.n19 bias1.t670 4.7605
R77 bias1.n19 bias1.t9 4.7605
R78 bias1.n19 bias1.t455 4.7605
R79 bias1.n19 bias1.t704 4.7605
R80 bias1.n19 bias1.t431 4.7605
R81 bias1.n20 bias1.t134 4.7605
R82 bias1.n20 bias1.t484 4.7605
R83 bias1.n20 bias1.t175 4.7605
R84 bias1.n20 bias1.t728 4.7605
R85 bias1.n20 bias1.t157 4.7605
R86 bias1.n20 bias1.t532 4.7605
R87 bias1.n20 bias1.t1122 4.7605
R88 bias1.n20 bias1.t571 4.7605
R89 bias1.n21 bias1.t1103 4.7605
R90 bias1.n21 bias1.t554 4.7605
R91 bias1.n21 bias1.t327 4.7605
R92 bias1.n21 bias1.t867 4.7605
R93 bias1.n21 bias1.t311 4.7605
R94 bias1.n21 bias1.t306 4.7605
R95 bias1.n21 bias1.t63 4.7605
R96 bias1.n21 bias1.t694 4.7605
R97 bias1.n8 bias1.t40 4.7605
R98 bias1.n8 bias1.t955 4.7605
R99 bias1.n8 bias1.t92 4.7605
R100 bias1.n8 bias1.t992 4.7605
R101 bias1.n8 bias1.t450 4.7605
R102 bias1.n8 bias1.t445 4.7605
R103 bias1.n32 bias1.t1111 4.65184
R104 bias1.n44 bias1.t265 4.65184
R105 bias1.n56 bias1.t19 4.65184
R106 bias1.n68 bias1.t369 4.65184
R107 bias1.n80 bias1.t1201 4.65184
R108 bias1.n92 bias1.t486 4.65184
R109 bias1.n104 bias1.t788 4.65184
R110 bias1.n116 bias1.t584 4.65184
R111 bias1.n128 bias1.t898 4.65184
R112 bias1.n140 bias1.t18 4.65184
R113 bias1.n22 bias1.t664 4.65134
R114 bias1.n22 bias1.t67 4.49693
R115 bias1.n22 bias1.t974 4.49693
R116 bias1.n22 bias1.t49 4.49693
R117 bias1.n22 bias1.t424 4.49693
R118 bias1.n22 bias1.t185 4.49693
R119 bias1.n22 bias1.t476 4.49693
R120 bias1.n23 bias1.t165 4.49693
R121 bias1.n23 bias1.t722 4.49693
R122 bias1.n23 bias1.t214 4.49693
R123 bias1.n23 bias1.t1116 4.49693
R124 bias1.n23 bias1.t506 4.49693
R125 bias1.n23 bias1.t564 4.49693
R126 bias1.n23 bias1.t1096 4.49693
R127 bias1.n23 bias1.t607 4.49693
R128 bias1.n24 bias1.t320 4.49693
R129 bias1.n24 bias1.t859 4.49693
R130 bias1.n24 bias1.t303 4.49693
R131 bias1.n24 bias1.t904 4.49693
R132 bias1.n24 bias1.t631 4.49693
R133 bias1.n24 bias1.t687 4.49693
R134 bias1.n24 bias1.t33 4.49693
R135 bias1.n24 bias1.t1003 4.49693
R136 bias1.n25 bias1.t83 4.49693
R137 bias1.n25 bias1.t985 4.49693
R138 bias1.n25 bias1.t441 4.49693
R139 bias1.n25 bias1.t1031 4.49693
R140 bias1.n25 bias1.t752 4.49693
R141 bias1.n25 bias1.t490 4.49693
R142 bias1.n25 bias1.t179 4.49693
R143 bias1.n25 bias1.t1084 4.49693
R144 bias1.n26 bias1.t236 4.49693
R145 bias1.n26 bias1.t1131 4.49693
R146 bias1.n26 bias1.t517 4.49693
R147 bias1.n26 bias1.t1112 4.49693
R148 bias1.n26 bias1.t893 4.49693
R149 bias1.n26 bias1.t891 4.49693
R150 bias1.n26 bias1.t333 4.49693
R151 bias1.n26 bias1.t873 4.49693
R152 bias1.n27 bias1.t374 4.49693
R153 bias1.n27 bias1.t70 4.49693
R154 bias1.n27 bias1.t642 4.49693
R155 bias1.n27 bias1.t50 4.49693
R156 bias1.n27 bias1.t679 4.49693
R157 bias1.n27 bias1.t1018 4.49693
R158 bias1.n27 bias1.t477 4.49693
R159 bias1.n27 bias1.t998 4.49693
R160 bias1.n28 bias1.t724 4.49693
R161 bias1.n28 bias1.t1043 4.49693
R162 bias1.n28 bias1.t764 4.49693
R163 bias1.n28 bias1.t197 4.49693
R164 bias1.n28 bias1.t746 4.49693
R165 bias1.n28 bias1.t1166 4.49693
R166 bias1.n28 bias1.t253 4.49693
R167 bias1.n28 bias1.t1144 4.49693
R168 bias1.n29 bias1.t861 4.49693
R169 bias1.n29 bias1.t1192 4.49693
R170 bias1.n29 bias1.t906 4.49693
R171 bias1.n29 bias1.t280 4.49693
R172 bias1.n29 bias1.t887 4.49693
R173 bias1.n29 bias1.t106 4.49693
R174 bias1.n29 bias1.t669 4.49693
R175 bias1.n29 bias1.t84 4.49693
R176 bias1.n30 bias1.t653 4.49693
R177 bias1.n30 bias1.t131 4.49693
R178 bias1.n30 bias1.t1036 4.49693
R179 bias1.n30 bias1.t416 4.49693
R180 bias1.n30 bias1.t1014 4.49693
R181 bias1.n30 bias1.t397 4.49693
R182 bias1.n30 bias1.t470 4.49693
R183 bias1.n30 bias1.t1066 4.49693
R184 bias1.n31 bias1.t447 4.49693
R185 bias1.n31 bias1.t145 4.49693
R186 bias1.n31 bias1.t500 4.49693
R187 bias1.n31 bias1.t192 4.49693
R188 bias1.n31 bias1.t807 4.49693
R189 bias1.n31 bias1.t171 4.49693
R190 bias1.n31 bias1.t603 4.49693
R191 bias1.n31 bias1.t850 4.49693
R192 bias1.t57 bias1.t587 4.49693
R193 bias1.t57 bias1.t297 4.49693
R194 bias1.t57 bias1.t626 4.49693
R195 bias1.t57 bias1.t344 4.49693
R196 bias1.t57 bias1.t880 4.49693
R197 bias1.n32 bias1.t123 4.49693
R198 bias1.n32 bias1.t685 4.49693
R199 bias1.n32 bias1.t110 4.49693
R200 bias1.n33 bias1.t104 4.49693
R201 bias1.n33 bias1.t1069 4.49693
R202 bias1.n33 bias1.t528 4.49693
R203 bias1.n33 bias1.t1049 4.49693
R204 bias1.n33 bias1.t771 4.49693
R205 bias1.n33 bias1.t1093 4.49693
R206 bias1.n33 bias1.t813 4.49693
R207 bias1.n33 bias1.t262 4.49693
R208 bias1.n34 bias1.t258 4.49693
R209 bias1.n34 bias1.t1151 4.49693
R210 bias1.n34 bias1.t298 4.49693
R211 bias1.n34 bias1.t1202 4.49693
R212 bias1.n34 bias1.t911 4.49693
R213 bias1.n34 bias1.t1181 4.49693
R214 bias1.n34 bias1.t947 4.49693
R215 bias1.n34 bias1.t329 4.49693
R216 bias1.n35 bias1.t392 4.49693
R217 bias1.n35 bias1.t93 4.49693
R218 bias1.n35 bias1.t710 4.49693
R219 bias1.n35 bias1.t139 4.49693
R220 bias1.n35 bias1.t695 4.49693
R221 bias1.n35 bias1.t119 4.49693
R222 bias1.n35 bias1.t1082 4.49693
R223 bias1.n35 bias1.t473 4.49693
R224 bias1.n36 bias1.t536 4.49693
R225 bias1.n36 bias1.t1062 4.49693
R226 bias1.n36 bias1.t785 4.49693
R227 bias1.n36 bias1.t291 4.49693
R228 bias1.n36 bias1.t825 4.49693
R229 bias1.n36 bias1.t563 4.49693
R230 bias1.n36 bias1.t805 4.49693
R231 bias1.n36 bias1.t604 4.49693
R232 bias1.n37 bias1.t663 4.49693
R233 bias1.n37 bias1.t1212 4.49693
R234 bias1.n37 bias1.t926 4.49693
R235 bias1.n37 bias1.t45 4.49693
R236 bias1.n37 bias1.t960 4.49693
R237 bias1.n37 bias1.t686 4.49693
R238 bias1.n37 bias1.t945 4.49693
R239 bias1.n37 bias1.t723 4.49693
R240 bias1.n38 bias1.t721 4.49693
R241 bias1.n38 bias1.t147 4.49693
R242 bias1.n38 bias1.t1052 4.49693
R243 bias1.n38 bias1.t436 4.49693
R244 bias1.n38 bias1.t1100 4.49693
R245 bias1.n38 bias1.t487 4.49693
R246 bias1.n38 bias1.t1080 4.49693
R247 bias1.n38 bias1.t801 4.49693
R248 bias1.n39 bias1.t858 4.49693
R249 bias1.n39 bias1.t301 4.49693
R250 bias1.n39 bias1.t838 4.49693
R251 bias1.n39 bias1.t574 4.49693
R252 bias1.n39 bias1.t34 4.49693
R253 bias1.n39 bias1.t616 4.49693
R254 bias1.n39 bias1.t331 4.49693
R255 bias1.n39 bias1.t597 4.49693
R256 bias1.n40 bias1.t984 4.49693
R257 bias1.n40 bias1.t440 4.49693
R258 bias1.n40 bias1.t969 4.49693
R259 bias1.n40 bias1.t699 4.49693
R260 bias1.n40 bias1.t1012 4.49693
R261 bias1.n40 bias1.t733 4.49693
R262 bias1.n40 bias1.t475 4.49693
R263 bias1.n40 bias1.t718 4.49693
R264 bias1.n41 bias1.t454 4.49693
R265 bias1.n41 bias1.t266 4.49693
R266 bias1.n41 bias1.t874 4.49693
R267 bias1.n41 bias1.t606 4.49693
R268 bias1.n41 bias1.t1141 4.49693
R269 bias1.n41 bias1.t644 4.49693
R270 bias1.n41 bias1.t1188 4.49693
R271 bias1.n41 bias1.t628 4.49693
R272 bias1.n42 bias1.t347 4.49693
R273 bias1.n42 bias1.t400 4.49693
R274 bias1.n42 bias1.t1000 4.49693
R275 bias1.n42 bias1.t385 4.49693
R276 bias1.n42 bias1.t82 4.49693
R277 bias1.n42 bias1.t766 4.49693
R278 bias1.n42 bias1.t127 4.49693
R279 bias1.n42 bias1.t1030 4.49693
R280 bias1.n43 bias1.t113 4.49693
R281 bias1.n43 bias1.t489 4.49693
R282 bias1.n43 bias1.t1147 4.49693
R283 bias1.n43 bias1.t529 4.49693
R284 bias1.n43 bias1.t235 4.49693
R285 bias1.n43 bias1.t516 4.49693
R286 bias1.n43 bias1.t282 4.49693
R287 bias1.n43 bias1.t1177 4.49693
R288 bias1.n7 bias1.t264 4.49693
R289 bias1.n7 bias1.t619 4.49693
R290 bias1.n7 bias1.t10 4.49693
R291 bias1.n7 bias1.t655 4.49693
R292 bias1.n7 bias1.t373 4.49693
R293 bias1.n7 bias1.t914 4.49693
R294 bias1.n7 bias1.t418 4.49693
R295 bias1.n7 bias1.t949 4.49693
R296 bias1.n7 bias1.t399 4.49693
R297 bias1.n7 bias1.t735 4.49693
R298 bias1.n44 bias1.t474 4.49693
R299 bias1.n44 bias1.t994 4.49693
R300 bias1.n44 bias1.t453 4.49693
R301 bias1.n45 bias1.t451 4.49693
R302 bias1.n45 bias1.t212 4.49693
R303 bias1.n45 bias1.t828 4.49693
R304 bias1.n45 bias1.t193 4.49693
R305 bias1.n45 bias1.t1094 4.49693
R306 bias1.n45 bias1.t248 4.49693
R307 bias1.n45 bias1.t1140 4.49693
R308 bias1.n45 bias1.t590 4.49693
R309 bias1.n46 bias1.t588 4.49693
R310 bias1.n46 bias1.t299 4.49693
R311 bias1.n46 bias1.t627 4.49693
R312 bias1.n46 bias1.t345 4.49693
R313 bias1.n46 bias1.t31 4.49693
R314 bias1.n46 bias1.t324 4.49693
R315 bias1.n46 bias1.t81 4.49693
R316 bias1.n46 bias1.t651 4.49693
R317 bias1.n47 bias1.t708 4.49693
R318 bias1.n47 bias1.t439 4.49693
R319 bias1.n47 bias1.t1028 4.49693
R320 bias1.n47 bias1.t488 4.49693
R321 bias1.n47 bias1.t1010 4.49693
R322 bias1.n47 bias1.t468 4.49693
R323 bias1.n47 bias1.t234 4.49693
R324 bias1.n47 bias1.t774 4.49693
R325 bias1.n48 bias1.t842 4.49693
R326 bias1.n48 bias1.t210 4.49693
R327 bias1.n48 bias1.t1109 4.49693
R328 bias1.n48 bias1.t618 4.49693
R329 bias1.n48 bias1.t1159 4.49693
R330 bias1.n48 bias1.t872 4.49693
R331 bias1.n48 bias1.t1136 4.49693
R332 bias1.n48 bias1.t913 4.49693
R333 bias1.n49 bias1.t971 4.49693
R334 bias1.n49 bias1.t355 4.49693
R335 bias1.n49 bias1.t48 4.49693
R336 bias1.n49 bias1.t396 4.49693
R337 bias1.n49 bias1.t99 4.49693
R338 bias1.n49 bias1.t997 4.49693
R339 bias1.n49 bias1.t78 4.49693
R340 bias1.n49 bias1.t1042 4.49693
R341 bias1.n50 bias1.t1040 4.49693
R342 bias1.n50 bias1.t502 4.49693
R343 bias1.n50 bias1.t196 4.49693
R344 bias1.n50 bias1.t742 4.49693
R345 bias1.n50 bias1.t252 4.49693
R346 bias1.n50 bias1.t789 4.49693
R347 bias1.n50 bias1.t229 4.49693
R348 bias1.n50 bias1.t1128 4.49693
R349 bias1.n51 bias1.t1190 4.49693
R350 bias1.n51 bias1.t630 4.49693
R351 bias1.n51 bias1.t1173 4.49693
R352 bias1.n51 bias1.t884 4.49693
R353 bias1.n51 bias1.t387 4.49693
R354 bias1.n51 bias1.t929 4.49693
R355 bias1.n51 bias1.t652 4.49693
R356 bias1.n51 bias1.t910 4.49693
R357 bias1.n52 bias1.t126 4.49693
R358 bias1.n52 bias1.t749 4.49693
R359 bias1.n52 bias1.t112 4.49693
R360 bias1.n52 bias1.t1013 4.49693
R361 bias1.n52 bias1.t151 4.49693
R362 bias1.n52 bias1.t1054 4.49693
R363 bias1.n52 bias1.t775 4.49693
R364 bias1.n52 bias1.t1039 4.49693
R365 bias1.n53 bias1.t761 4.49693
R366 bias1.n53 bias1.t138 4.49693
R367 bias1.n53 bias1.t757 4.49693
R368 bias1.n53 bias1.t499 4.49693
R369 bias1.n53 bias1.t1019 4.49693
R370 bias1.n53 bias1.t537 4.49693
R371 bias1.n53 bias1.t1064 4.49693
R372 bias1.n53 bias1.t522 4.49693
R373 bias1.n54 bias1.t224 4.49693
R374 bias1.n54 bias1.t290 4.49693
R375 bias1.n54 bias1.t899 4.49693
R376 bias1.n54 bias1.t272 4.49693
R377 bias1.n54 bias1.t1169 4.49693
R378 bias1.n54 bias1.t662 4.49693
R379 bias1.n54 bias1.t1213 4.49693
R380 bias1.n54 bias1.t925 4.49693
R381 bias1.n55 bias1.t1195 4.49693
R382 bias1.n55 bias1.t362 4.49693
R383 bias1.n55 bias1.t1025 4.49693
R384 bias1.n55 bias1.t408 4.49693
R385 bias1.n55 bias1.t111 4.49693
R386 bias1.n55 bias1.t390 4.49693
R387 bias1.n55 bias1.t148 4.49693
R388 bias1.n55 bias1.t1053 4.49693
R389 bias1.n6 bias1.t136 4.49693
R390 bias1.n6 bias1.t512 4.49693
R391 bias1.n6 bias1.t1095 4.49693
R392 bias1.n6 bias1.t547 4.49693
R393 bias1.n6 bias1.t263 4.49693
R394 bias1.n6 bias1.t796 4.49693
R395 bias1.n6 bias1.t302 4.49693
R396 bias1.n6 bias1.t837 4.49693
R397 bias1.n7 bias1.t288 4.49693
R398 bias1.n7 bias1.t638 4.49693
R399 bias1.n56 bias1.t247 4.49693
R400 bias1.n56 bias1.t782 4.49693
R401 bias1.n56 bias1.t222 4.49693
R402 bias1.n57 bias1.t216 4.49693
R403 bias1.n57 bias1.t1186 4.49693
R404 bias1.n57 bias1.t625 4.49693
R405 bias1.n57 bias1.t1167 4.49693
R406 bias1.n57 bias1.t877 4.49693
R407 bias1.n57 bias1.t1209 4.49693
R408 bias1.n57 bias1.t922 4.49693
R409 bias1.n57 bias1.t364 4.49693
R410 bias1.n58 bias1.t360 4.49693
R411 bias1.n58 bias1.t54 4.49693
R412 bias1.n58 bias1.t403 4.49693
R413 bias1.n58 bias1.t107 4.49693
R414 bias1.n58 bias1.t1006 4.49693
R415 bias1.n58 bias1.t86 4.49693
R416 bias1.n58 bias1.t1050 4.49693
R417 bias1.n58 bias1.t433 4.49693
R418 bias1.n59 bias1.t509 4.49693
R419 bias1.n59 bias1.t204 4.49693
R420 bias1.n59 bias1.t812 4.49693
R421 bias1.n59 bias1.t260 4.49693
R422 bias1.n59 bias1.t794 4.49693
R423 bias1.n59 bias1.t240 4.49693
R424 bias1.n59 bias1.t1203 4.49693
R425 bias1.n59 bias1.t573 4.49693
R426 bias1.n60 bias1.t636 4.49693
R427 bias1.n60 bias1.t1178 4.49693
R428 bias1.n60 bias1.t895 4.49693
R429 bias1.n60 bias1.t394 4.49693
R430 bias1.n60 bias1.t935 4.49693
R431 bias1.n60 bias1.t660 4.49693
R432 bias1.n60 bias1.t917 4.49693
R433 bias1.n60 bias1.t696 4.49693
R434 bias1.n61 bias1.t759 4.49693
R435 bias1.n61 bias1.t117 4.49693
R436 bias1.n61 bias1.t1021 4.49693
R437 bias1.n61 bias1.t160 4.49693
R438 bias1.n61 bias1.t1065 4.49693
R439 bias1.n61 bias1.t786 4.49693
R440 bias1.n61 bias1.t1046 4.49693
R441 bias1.n61 bias1.t826 4.49693
R442 bias1.n62 bias1.t823 4.49693
R443 bias1.n62 bias1.t273 4.49693
R444 bias1.n62 bias1.t1170 4.49693
R445 bias1.n62 bias1.t543 4.49693
R446 bias1.n62 bias1.t1214 4.49693
R447 bias1.n62 bias1.t586 4.49693
R448 bias1.n62 bias1.t1199 4.49693
R449 bias1.n62 bias1.t909 4.49693
R450 bias1.n63 bias1.t959 4.49693
R451 bias1.n63 bias1.t409 4.49693
R452 bias1.n63 bias1.t944 4.49693
R453 bias1.n63 bias1.t672 4.49693
R454 bias1.n63 bias1.t149 4.49693
R455 bias1.n63 bias1.t707 4.49693
R456 bias1.n63 bias1.t438 4.49693
R457 bias1.n63 bias1.t688 4.49693
R458 bias1.n64 bias1.t1099 4.49693
R459 bias1.n64 bias1.t549 4.49693
R460 bias1.n64 bias1.t1078 4.49693
R461 bias1.n64 bias1.t799 4.49693
R462 bias1.n64 bias1.t1124 4.49693
R463 bias1.n64 bias1.t840 4.49693
R464 bias1.n64 bias1.t577 4.49693
R465 bias1.n64 bias1.t820 4.49693
R466 bias1.n65 bias1.t560 4.49693
R467 bias1.n65 bias1.t232 4.49693
R468 bias1.n65 bias1.t841 4.49693
R469 bias1.n65 bias1.t578 4.49693
R470 bias1.n65 bias1.t1108 4.49693
R471 bias1.n65 bias1.t617 4.49693
R472 bias1.n65 bias1.t1158 4.49693
R473 bias1.n65 bias1.t601 4.49693
R474 bias1.n66 bias1.t317 4.49693
R475 bias1.n66 bias1.t371 4.49693
R476 bias1.n66 bias1.t970 4.49693
R477 bias1.n66 bias1.t354 4.49693
R478 bias1.n66 bias1.t47 4.49693
R479 bias1.n66 bias1.t734 4.49693
R480 bias1.n66 bias1.t98 4.49693
R481 bias1.n66 bias1.t996 4.49693
R482 bias1.n67 bias1.t77 4.49693
R483 bias1.n67 bias1.t457 4.49693
R484 bias1.n67 bias1.t1113 4.49693
R485 bias1.n67 bias1.t501 4.49693
R486 bias1.n67 bias1.t195 4.49693
R487 bias1.n67 bias1.t485 4.49693
R488 bias1.n67 bias1.t251 4.49693
R489 bias1.n67 bias1.t1143 4.49693
R490 bias1.n0 bias1.t230 4.49693
R491 bias1.n0 bias1.t591 4.49693
R492 bias1.n0 bias1.t1189 4.49693
R493 bias1.n0 bias1.t629 4.49693
R494 bias1.n0 bias1.t348 4.49693
R495 bias1.n0 bias1.t883 4.49693
R496 bias1.n0 bias1.t386 4.49693
R497 bias1.n0 bias1.t928 4.49693
R498 bias1.n1 bias1.t370 4.49693
R499 bias1.n1 bias1.t712 4.49693
R500 bias1.n68 bias1.t576 4.49693
R501 bias1.n68 bias1.t1107 4.49693
R502 bias1.n68 bias1.t559 4.49693
R503 bias1.n69 bias1.t556 4.49693
R504 bias1.n69 bias1.t330 4.49693
R505 bias1.n69 bias1.t938 4.49693
R506 bias1.n69 bias1.t312 4.49693
R507 bias1.n69 bias1.t1211 4.49693
R508 bias1.n69 bias1.t352 4.49693
R509 bias1.n69 bias1.t44 4.49693
R510 bias1.n69 bias1.t684 4.49693
R511 bias1.n70 bias1.t681 4.49693
R512 bias1.n70 bias1.t405 4.49693
R513 bias1.n70 bias1.t716 4.49693
R514 bias1.n70 bias1.t452 4.49693
R515 bias1.n70 bias1.t146 4.49693
R516 bias1.n70 bias1.t429 4.49693
R517 bias1.n70 bias1.t194 4.49693
R518 bias1.n70 bias1.t741 4.49693
R519 bias1.n71 bias1.t808 4.49693
R520 bias1.n71 bias1.t545 4.49693
R521 bias1.n71 bias1.t1139 4.49693
R522 bias1.n71 bias1.t589 4.49693
R523 bias1.n71 bias1.t1120 4.49693
R524 bias1.n71 bias1.t568 4.49693
R525 bias1.n71 bias1.t346 4.49693
R526 bias1.n71 bias1.t882 4.49693
R527 bias1.n72 bias1.t946 4.49693
R528 bias1.n72 bias1.t323 4.49693
R529 bias1.n72 bias1.t15 4.49693
R530 bias1.n72 bias1.t709 4.49693
R531 bias1.n72 bias1.t61 4.49693
R532 bias1.n72 bias1.t968 4.49693
R533 bias1.n72 bias1.t38 4.49693
R534 bias1.n72 bias1.t1011 4.49693
R535 bias1.n73 bias1.t1081 4.49693
R536 bias1.n73 bias1.t467 4.49693
R537 bias1.n73 bias1.t162 4.49693
R538 bias1.n73 bias1.t515 4.49693
R539 bias1.n73 bias1.t211 4.49693
R540 bias1.n73 bias1.t1110 4.49693
R541 bias1.n73 bias1.t188 4.49693
R542 bias1.n73 bias1.t1160 4.49693
R543 bias1.n74 bias1.t1157 4.49693
R544 bias1.n74 bias1.t600 4.49693
R545 bias1.n74 bias1.t316 4.49693
R546 bias1.n74 bias1.t849 4.49693
R547 bias1.n74 bias1.t357 4.49693
R548 bias1.n74 bias1.t900 4.49693
R549 bias1.n74 bias1.t340 4.49693
R550 bias1.n74 bias1.t28 4.49693
R551 bias1.n75 bias1.t96 4.49693
R552 bias1.n75 bias1.t720 4.49693
R553 bias1.n75 bias1.t74 4.49693
R554 bias1.n75 bias1.t980 4.49693
R555 bias1.n75 bias1.t504 4.49693
R556 bias1.n75 bias1.t1026 4.49693
R557 bias1.n75 bias1.t744 4.49693
R558 bias1.n75 bias1.t1005 4.49693
R559 bias1.n76 bias1.t250 4.49693
R560 bias1.n76 bias1.t857 4.49693
R561 bias1.n76 bias1.t227 4.49693
R562 bias1.n76 bias1.t1126 4.49693
R563 bias1.n76 bias1.t277 4.49693
R564 bias1.n76 bias1.t1174 4.49693
R565 bias1.n76 bias1.t885 4.49693
R566 bias1.n76 bias1.t1154 4.49693
R567 bias1.n77 bias1.t870 4.49693
R568 bias1.n77 bias1.t105 4.49693
R569 bias1.n77 bias1.t727 4.49693
R570 bias1.n77 bias1.t463 4.49693
R571 bias1.n77 bias1.t986 4.49693
R572 bias1.n77 bias1.t511 4.49693
R573 bias1.n77 bias1.t1035 4.49693
R574 bias1.n77 bias1.t492 4.49693
R575 bias1.n78 bias1.t184 4.49693
R576 bias1.n78 bias1.t259 4.49693
R577 bias1.n78 bias1.t865 4.49693
R578 bias1.n78 bias1.t238 4.49693
R579 bias1.n78 bias1.t1133 4.49693
R580 bias1.n78 bias1.t637 4.49693
R581 bias1.n78 bias1.t1182 4.49693
R582 bias1.n78 bias1.t897 4.49693
R583 bias1.n79 bias1.t1161 4.49693
R584 bias1.n79 bias1.t335 4.49693
R585 bias1.n79 bias1.t990 4.49693
R586 bias1.n79 bias1.t379 4.49693
R587 bias1.n79 bias1.t73 4.49693
R588 bias1.n79 bias1.t358 4.49693
R589 bias1.n79 bias1.t120 4.49693
R590 bias1.n79 bias1.t1024 4.49693
R591 bias1.n9 bias1.t101 4.49693
R592 bias1.n9 bias1.t481 4.49693
R593 bias1.n9 bias1.t1063 4.49693
R594 bias1.n9 bias1.t523 4.49693
R595 bias1.n9 bias1.t225 4.49693
R596 bias1.n9 bias1.t767 4.49693
R597 bias1.n9 bias1.t275 4.49693
R598 bias1.n9 bias1.t806 4.49693
R599 bias1.n1 bias1.t256 4.49693
R600 bias1.n1 bias1.t612 4.49693
R601 bias1.n80 bias1.t206 4.49693
R602 bias1.n80 bias1.t753 4.49693
R603 bias1.n80 bias1.t183 4.49693
R604 bias1.n81 bias1.t181 4.49693
R605 bias1.n81 bias1.t1152 4.49693
R606 bias1.n81 bias1.t596 4.49693
R607 bias1.n81 bias1.t1132 4.49693
R608 bias1.n81 bias1.t847 4.49693
R609 bias1.n81 bias1.t1180 4.49693
R610 bias1.n81 bias1.t896 4.49693
R611 bias1.n81 bias1.t336 4.49693
R612 bias1.n82 bias1.t334 4.49693
R613 bias1.n82 bias1.t23 4.49693
R614 bias1.n82 bias1.t377 4.49693
R615 bias1.n82 bias1.t72 4.49693
R616 bias1.n82 bias1.t978 4.49693
R617 bias1.n82 bias1.t51 4.49693
R618 bias1.n82 bias1.t1023 4.49693
R619 bias1.n82 bias1.t402 4.49693
R620 bias1.n83 bias1.t478 4.49693
R621 bias1.n83 bias1.t170 4.49693
R622 bias1.n83 bias1.t784 4.49693
R623 bias1.n83 bias1.t223 4.49693
R624 bias1.n83 bias1.t765 4.49693
R625 bias1.n83 bias1.t200 4.49693
R626 bias1.n83 bias1.t1172 4.49693
R627 bias1.n83 bias1.t544 4.49693
R628 bias1.n84 bias1.t609 4.49693
R629 bias1.n84 bias1.t1146 4.49693
R630 bias1.n84 bias1.t862 4.49693
R631 bias1.n84 bias1.t366 4.49693
R632 bias1.n84 bias1.t907 4.49693
R633 bias1.n84 bias1.t634 4.49693
R634 bias1.n84 bias1.t890 4.49693
R635 bias1.n84 bias1.t673 4.49693
R636 bias1.n85 bias1.t730 4.49693
R637 bias1.n85 bias1.t87 4.49693
R638 bias1.n85 bias1.t987 4.49693
R639 bias1.n85 bias1.t135 4.49693
R640 bias1.n85 bias1.t1038 4.49693
R641 bias1.n85 bias1.t756 4.49693
R642 bias1.n85 bias1.t1017 4.49693
R643 bias1.n85 bias1.t800 4.49693
R644 bias1.n86 bias1.t795 4.49693
R645 bias1.n86 bias1.t241 4.49693
R646 bias1.n86 bias1.t1134 4.49693
R647 bias1.n86 bias1.t520 4.49693
R648 bias1.n86 bias1.t1184 4.49693
R649 bias1.n86 bias1.t558 4.49693
R650 bias1.n86 bias1.t1165 4.49693
R651 bias1.n86 bias1.t875 4.49693
R652 bias1.n87 bias1.t937 4.49693
R653 bias1.n87 bias1.t381 4.49693
R654 bias1.n87 bias1.t918 4.49693
R655 bias1.n87 bias1.t647 4.49693
R656 bias1.n87 bias1.t122 4.49693
R657 bias1.n87 bias1.t683 4.49693
R658 bias1.n87 bias1.t407 4.49693
R659 bias1.n87 bias1.t668 4.49693
R660 bias1.n88 bias1.t1068 4.49693
R661 bias1.n88 bias1.t526 4.49693
R662 bias1.n88 bias1.t1047 4.49693
R663 bias1.n88 bias1.t769 4.49693
R664 bias1.n88 bias1.t1092 4.49693
R665 bias1.n88 bias1.t809 4.49693
R666 bias1.n88 bias1.t546 4.49693
R667 bias1.n88 bias1.t792 4.49693
R668 bias1.n89 bias1.t533 4.49693
R669 bias1.n89 bias1.t705 4.49693
R670 bias1.n89 bias1.t130 4.49693
R671 bias1.n89 bias1.t1033 4.49693
R672 bias1.n89 bias1.t415 4.49693
R673 bias1.n89 bias1.t1076 4.49693
R674 bias1.n89 bias1.t462 4.49693
R675 bias1.n89 bias1.t1057 4.49693
R676 bias1.n90 bias1.t776 4.49693
R677 bias1.n90 bias1.t836 4.49693
R678 bias1.n90 bias1.t285 4.49693
R679 bias1.n90 bias1.t815 4.49693
R680 bias1.n90 bias1.t553 4.49693
R681 bias1.n90 bias1.t16 4.49693
R682 bias1.n90 bias1.t595 4.49693
R683 bias1.n90 bias1.t310 4.49693
R684 bias1.n91 bias1.t580 4.49693
R685 bias1.n91 bias1.t915 4.49693
R686 bias1.n91 bias1.t421 4.49693
R687 bias1.n91 bias1.t951 4.49693
R688 bias1.n91 bias1.t680 4.49693
R689 bias1.n91 bias1.t940 4.49693
R690 bias1.n91 bias1.t715 4.49693
R691 bias1.n91 bias1.t449 4.49693
R692 bias1.n1 bias1.t701 4.49693
R693 bias1.n1 bias1.t1044 4.49693
R694 bias1.n1 bias1.t497 4.49693
R695 bias1.n1 bias1.t1087 4.49693
R696 bias1.n1 bias1.t804 4.49693
R697 bias1.n1 bias1.t168 4.49693
R698 bias1.n1 bias1.t853 4.49693
R699 bias1.n1 bias1.t221 4.49693
R700 bias1.n1 bias1.t833 4.49693
R701 bias1.n1 bias1.t1194 4.49693
R702 bias1.n92 bias1.t674 4.49693
R703 bias1.n92 bias1.t13 4.49693
R704 bias1.n92 bias1.t658 4.49693
R705 bias1.n93 bias1.t656 4.49693
R706 bias1.n93 bias1.t435 4.49693
R707 bias1.n93 bias1.t1037 4.49693
R708 bias1.n93 bias1.t419 4.49693
R709 bias1.n93 bias1.t116 4.49693
R710 bias1.n93 bias1.t465 4.49693
R711 bias1.n93 bias1.t159 4.49693
R712 bias1.n93 bias1.t781 4.49693
R713 bias1.n94 bias1.t778 4.49693
R714 bias1.n94 bias1.t519 4.49693
R715 bias1.n94 bias1.t818 4.49693
R716 bias1.n94 bias1.t557 4.49693
R717 bias1.n94 bias1.t271 4.49693
R718 bias1.n94 bias1.t540 4.49693
R719 bias1.n94 bias1.t314 4.49693
R720 bias1.n94 bias1.t848 4.49693
R721 bias1.n95 bias1.t919 4.49693
R722 bias1.n95 bias1.t646 4.49693
R723 bias1.n95 bias1.t43 4.49693
R724 bias1.n95 bias1.t682 4.49693
R725 bias1.n95 bias1.t24 4.49693
R726 bias1.n95 bias1.t667 4.49693
R727 bias1.n95 bias1.t456 4.49693
R728 bias1.n95 bias1.t979 4.49693
R729 bias1.n96 bias1.t1048 4.49693
R730 bias1.n96 bias1.t428 4.49693
R731 bias1.n96 bias1.t132 4.49693
R732 bias1.n96 bias1.t810 4.49693
R733 bias1.n96 bias1.t173 4.49693
R734 bias1.n96 bias1.t1077 4.49693
R735 bias1.n96 bias1.t155 4.49693
R736 bias1.n96 bias1.t1123 4.49693
R737 bias1.n97 bias1.t1200 4.49693
R738 bias1.n97 bias1.t567 4.49693
R739 bias1.n97 bias1.t286 4.49693
R740 bias1.n97 bias1.t615 4.49693
R741 bias1.n97 bias1.t325 4.49693
R742 bias1.n97 bias1.t17 4.49693
R743 bias1.n97 bias1.t307 4.49693
R744 bias1.n97 bias1.t64 4.49693
R745 bias1.n98 bias1.t60 4.49693
R746 bias1.n98 bias1.t691 4.49693
R747 bias1.n98 bias1.t422 4.49693
R748 bias1.n98 bias1.t952 4.49693
R749 bias1.n98 bias1.t469 4.49693
R750 bias1.n98 bias1.t989 4.49693
R751 bias1.n98 bias1.t446 4.49693
R752 bias1.n98 bias1.t143 4.49693
R753 bias1.n99 bias1.t209 4.49693
R754 bias1.n99 bias1.t821 4.49693
R755 bias1.n99 bias1.t187 4.49693
R756 bias1.n99 bias1.t1088 4.49693
R757 bias1.n99 bias1.t602 4.49693
R758 bias1.n99 bias1.t1135 4.49693
R759 bias1.n99 bias1.t854 4.49693
R760 bias1.n99 bias1.t1117 4.49693
R761 bias1.n100 bias1.t353 4.49693
R762 bias1.n100 bias1.t957 4.49693
R763 bias1.n100 bias1.t339 4.49693
R764 bias1.n100 bias1.t27 4.49693
R765 bias1.n100 bias1.t384 4.49693
R766 bias1.n100 bias1.t76 4.49693
R767 bias1.n100 bias1.t983 4.49693
R768 bias1.n100 bias1.t56 4.49693
R769 bias1.n101 bias1.t967 4.49693
R770 bias1.n101 bias1.t71 4.49693
R771 bias1.n101 bias1.t700 4.49693
R772 bias1.n101 bias1.t427 4.49693
R773 bias1.n101 bias1.t961 4.49693
R774 bias1.n101 bias1.t480 4.49693
R775 bias1.n101 bias1.t1001 4.49693
R776 bias1.n101 bias1.t459 4.49693
R777 bias1.n102 bias1.t153 4.49693
R778 bias1.n102 bias1.t218 4.49693
R779 bias1.n102 bias1.t832 4.49693
R780 bias1.n102 bias1.t198 4.49693
R781 bias1.n102 bias1.t1101 4.49693
R782 bias1.n102 bias1.t611 4.49693
R783 bias1.n102 bias1.t1148 4.49693
R784 bias1.n102 bias1.t863 4.49693
R785 bias1.n103 bias1.t1130 4.49693
R786 bias1.n103 bias1.t304 4.49693
R787 bias1.n103 bias1.t964 4.49693
R788 bias1.n103 bias1.t349 4.49693
R789 bias1.n103 bias1.t36 4.49693
R790 bias1.n103 bias1.t332 4.49693
R791 bias1.n103 bias1.t88 4.49693
R792 bias1.n103 bias1.t988 4.49693
R793 bias1.n3 bias1.t68 4.49693
R794 bias1.n3 bias1.t443 4.49693
R795 bias1.n3 bias1.t1034 4.49693
R796 bias1.n3 bias1.t494 4.49693
R797 bias1.n3 bias1.t186 4.49693
R798 bias1.n3 bias1.t736 4.49693
R799 bias1.n3 bias1.t243 4.49693
R800 bias1.n3 bias1.t779 4.49693
R801 bias1.n4 bias1.t215 4.49693
R802 bias1.n4 bias1.t583 4.49693
R803 bias1.n104 bias1.t982 4.49693
R804 bias1.n104 bias1.t365 4.49693
R805 bias1.n104 bias1.t966 4.49693
R806 bias1.n105 bias1.t963 4.49693
R807 bias1.n105 bias1.t743 4.49693
R808 bias1.n105 bias1.t177 4.49693
R809 bias1.n105 bias1.t729 4.49693
R810 bias1.n105 bias1.t464 4.49693
R811 bias1.n105 bias1.t770 4.49693
R812 bias1.n105 bias1.t514 4.49693
R813 bias1.n105 bias1.t1106 4.49693
R814 bias1.n106 bias1.t1104 4.49693
R815 bias1.n106 bias1.t817 4.49693
R816 bias1.n106 bias1.t1150 4.49693
R817 bias1.n106 bias1.t868 4.49693
R818 bias1.n106 bias1.t598 4.49693
R819 bias1.n106 bias1.t846 4.49693
R820 bias1.n106 bias1.t640 4.49693
R821 bias1.n106 bias1.t1183 4.49693
R822 bias1.n107 bias1.t41 4.49693
R823 bias1.n107 bias1.t956 4.49693
R824 bias1.n107 bias1.t395 4.49693
R825 bias1.n107 bias1.t993 4.49693
R826 bias1.n107 bias1.t380 4.49693
R827 bias1.n107 bias1.t977 4.49693
R828 bias1.n107 bias1.t760 4.49693
R829 bias1.n107 bias1.t121 4.49693
R830 bias1.n108 bias1.t191 4.49693
R831 bias1.n108 bias1.t739 4.49693
R832 bias1.n108 bias1.t482 4.49693
R833 bias1.n108 bias1.t1138 4.49693
R834 bias1.n108 bias1.t525 4.49693
R835 bias1.n108 bias1.t226 4.49693
R836 bias1.n108 bias1.t508 4.49693
R837 bias1.n108 bias1.t276 4.49693
R838 bias1.n109 bias1.t343 4.49693
R839 bias1.n109 bias1.t879 4.49693
R840 bias1.n109 bias1.t614 4.49693
R841 bias1.n109 bias1.t924 4.49693
R842 bias1.n109 bias1.t650 4.49693
R843 bias1.n109 bias1.t367 4.49693
R844 bias1.n109 bias1.t633 4.49693
R845 bias1.n109 bias1.t412 4.49693
R846 bias1.n110 bias1.t411 4.49693
R847 bias1.n110 bias1.t1008 4.49693
R848 bias1.n110 bias1.t732 4.49693
R849 bias1.n110 bias1.t90 4.49693
R850 bias1.n110 bias1.t773 4.49693
R851 bias1.n110 bias1.t137 4.49693
R852 bias1.n110 bias1.t755 4.49693
R853 bias1.n110 bias1.t498 4.49693
R854 bias1.n111 bias1.t550 4.49693
R855 bias1.n111 bias1.t1155 4.49693
R856 bias1.n111 bias1.t534 4.49693
R857 bias1.n111 bias1.t244 4.49693
R858 bias1.n111 bias1.t912 4.49693
R859 bias1.n111 bias1.t289 4.49693
R860 bias1.n111 bias1.t1187 4.49693
R861 bias1.n111 bias1.t270 4.49693
R862 bias1.n112 bias1.t676 4.49693
R863 bias1.n112 bias1.t95 4.49693
R864 bias1.n112 bias1.t661 4.49693
R865 bias1.n112 bias1.t383 4.49693
R866 bias1.n112 bias1.t698 4.49693
R867 bias1.n112 bias1.t423 4.49693
R868 bias1.n112 bias1.t124 4.49693
R869 bias1.n112 bias1.t406 4.49693
R870 bias1.n113 bias1.t109 4.49693
R871 bias1.n113 bias1.t1156 4.49693
R872 bias1.n113 bias1.t599 4.49693
R873 bias1.n113 bias1.t315 4.49693
R874 bias1.n113 bias1.t852 4.49693
R875 bias1.n113 bias1.t356 4.49693
R876 bias1.n113 bias1.t902 4.49693
R877 bias1.n113 bias1.t341 4.49693
R878 bias1.n114 bias1.t29 4.49693
R879 bias1.n114 bias1.t97 4.49693
R880 bias1.n114 bias1.t719 4.49693
R881 bias1.n114 bias1.t75 4.49693
R882 bias1.n114 bias1.t981 4.49693
R883 bias1.n114 bias1.t503 4.49693
R884 bias1.n114 bias1.t1027 4.49693
R885 bias1.n114 bias1.t745 4.49693
R886 bias1.n115 bias1.t1004 4.49693
R887 bias1.n115 bias1.t176 4.49693
R888 bias1.n115 bias1.t856 4.49693
R889 bias1.n115 bias1.t228 4.49693
R890 bias1.n115 bias1.t1127 4.49693
R891 bias1.n115 bias1.t203 4.49693
R892 bias1.n115 bias1.t1175 4.49693
R893 bias1.n115 bias1.t886 4.49693
R894 bias1.n4 bias1.t1153 4.49693
R895 bias1.n4 bias1.t328 4.49693
R896 bias1.n4 bias1.t927 4.49693
R897 bias1.n4 bias1.t368 4.49693
R898 bias1.n4 bias1.t65 4.49693
R899 bias1.n4 bias1.t639 4.49693
R900 bias1.n4 bias1.t114 4.49693
R901 bias1.n4 bias1.t675 4.49693
R902 bias1.n4 bias1.t94 4.49693
R903 bias1.n4 bias1.t472 4.49693
R904 bias1.n116 bias1.t768 4.49693
R905 bias1.n116 bias1.t129 4.49693
R906 bias1.n116 bias1.t751 4.49693
R907 bias1.n117 bias1.t747 4.49693
R908 bias1.n117 bias1.t541 4.49693
R909 bias1.n117 bias1.t1149 4.49693
R910 bias1.n117 bias1.t530 4.49693
R911 bias1.n117 bias1.t237 4.49693
R912 bias1.n117 bias1.t565 4.49693
R913 bias1.n117 bias1.t284 4.49693
R914 bias1.n117 bias1.t892 4.49693
R915 bias1.n118 bias1.t888 4.49693
R916 bias1.n118 bias1.t621 4.49693
R917 bias1.n118 bias1.t931 4.49693
R918 bias1.n118 bias1.t657 4.49693
R919 bias1.n118 bias1.t376 4.49693
R920 bias1.n118 bias1.t641 4.49693
R921 bias1.n118 bias1.t420 4.49693
R922 bias1.n118 bias1.t950 4.49693
R923 bias1.n119 bias1.t1015 4.49693
R924 bias1.n119 bias1.t737 4.49693
R925 bias1.n119 bias1.t158 4.49693
R926 bias1.n119 bias1.t780 4.49693
R927 bias1.n119 bias1.t140 4.49693
R928 bias1.n119 bias1.t762 4.49693
R929 bias1.n119 bias1.t561 4.49693
R930 bias1.n119 bias1.t1086 4.49693
R931 bias1.n120 bias1.t1163 4.49693
R932 bias1.n120 bias1.t538 4.49693
R933 bias1.n120 bias1.t255 4.49693
R934 bias1.n120 bias1.t920 4.49693
R935 bias1.n120 bias1.t292 4.49693
R936 bias1.n120 bias1.t1193 4.49693
R937 bias1.n120 bias1.t279 4.49693
R938 bias1.n120 bias1.t25 4.49693
R939 bias1.n121 bias1.t103 4.49693
R940 bias1.n121 bias1.t666 4.49693
R941 bias1.n121 bias1.t389 4.49693
R942 bias1.n121 bias1.t702 4.49693
R943 bias1.n121 bias1.t430 4.49693
R944 bias1.n121 bias1.t133 4.49693
R945 bias1.n121 bias1.t414 4.49693
R946 bias1.n121 bias1.t174 4.49693
R947 bias1.n122 bias1.t172 4.49693
R948 bias1.n122 bias1.t791 4.49693
R949 bias1.n122 bias1.t531 4.49693
R950 bias1.n122 bias1.t1056 4.49693
R951 bias1.n122 bias1.t569 4.49693
R952 bias1.n122 bias1.t1102 4.49693
R953 bias1.n122 bias1.t552 4.49693
R954 bias1.n122 bias1.t268 4.49693
R955 bias1.n123 bias1.t322 4.49693
R956 bias1.n123 bias1.t934 4.49693
R957 bias1.n123 bias1.t305 4.49693
R958 bias1.n123 bias1.t1206 4.49693
R959 bias1.n123 bias1.t692 4.49693
R960 bias1.n123 bias1.t37 4.49693
R961 bias1.n123 bias1.t953 4.49693
R962 bias1.n123 bias1.t21 4.49693
R963 bias1.n124 bias1.t466 4.49693
R964 bias1.n124 bias1.t1061 4.49693
R965 bias1.n124 bias1.t444 4.49693
R966 bias1.n124 bias1.t141 4.49693
R967 bias1.n124 bias1.t495 4.49693
R968 bias1.n124 bias1.t189 4.49693
R969 bias1.n124 bias1.t1089 4.49693
R970 bias1.n124 bias1.t166 4.49693
R971 bias1.n125 bias1.t1073 4.49693
R972 bias1.n125 bias1.t35 4.49693
R973 bias1.n125 bias1.t677 4.49693
R974 bias1.n125 bias1.t398 4.49693
R975 bias1.n125 bias1.t939 4.49693
R976 bias1.n125 bias1.t442 4.49693
R977 bias1.n125 bias1.t972 4.49693
R978 bias1.n125 bias1.t425 4.49693
R979 bias1.n126 bias1.t125 4.49693
R980 bias1.n126 bias1.t182 4.49693
R981 bias1.n126 bias1.t802 4.49693
R982 bias1.n126 bias1.t163 4.49693
R983 bias1.n126 bias1.t1070 4.49693
R984 bias1.n126 bias1.t582 4.49693
R985 bias1.n126 bias1.t1114 4.49693
R986 bias1.n126 bias1.t830 4.49693
R987 bias1.n127 bias1.t1098 4.49693
R988 bias1.n127 bias1.t278 4.49693
R989 bias1.n127 bias1.t941 4.49693
R990 bias1.n127 bias1.t318 4.49693
R991 bias1.n127 bias1.t7 4.49693
R992 bias1.n127 bias1.t300 4.49693
R993 bias1.n127 bias1.t52 4.49693
R994 bias1.n127 bias1.t962 4.49693
R995 bias1.n5 bias1.t32 4.49693
R996 bias1.n5 bias1.t413 4.49693
R997 bias1.n5 bias1.t1002 4.49693
R998 bias1.n5 bias1.t460 4.49693
R999 bias1.n5 bias1.t154 4.49693
R1000 bias1.n5 bias1.t713 4.49693
R1001 bias1.n5 bias1.t201 4.49693
R1002 bias1.n5 bias1.t750 4.49693
R1003 bias1.n2 bias1.t180 4.49693
R1004 bias1.n2 bias1.t551 4.49693
R1005 bias1.n128 bias1.t1090 4.49693
R1006 bias1.n128 bias1.t479 4.49693
R1007 bias1.n128 bias1.t1074 4.49693
R1008 bias1.n129 bias1.t1071 4.49693
R1009 bias1.n129 bias1.t851 4.49693
R1010 bias1.n129 bias1.t294 4.49693
R1011 bias1.n129 bias1.t831 4.49693
R1012 bias1.n129 bias1.t566 4.49693
R1013 bias1.n129 bias1.t876 4.49693
R1014 bias1.n129 bias1.t610 4.49693
R1015 bias1.n129 bias1.t12 4.49693
R1016 bias1.n130 bias1.t8 4.49693
R1017 bias1.n130 bias1.t932 4.49693
R1018 bias1.n130 bias1.t53 4.49693
R1019 bias1.n130 bias1.t965 4.49693
R1020 bias1.n130 bias1.t689 4.49693
R1021 bias1.n130 bias1.t948 4.49693
R1022 bias1.n130 bias1.t731 4.49693
R1023 bias1.n130 bias1.t89 4.49693
R1024 bias1.n131 bias1.t156 4.49693
R1025 bias1.n131 bias1.t1059 4.49693
R1026 bias1.n131 bias1.t513 4.49693
R1027 bias1.n131 bias1.t1105 4.49693
R1028 bias1.n131 bias1.t493 4.49693
R1029 bias1.n131 bias1.t1085 4.49693
R1030 bias1.n131 bias1.t869 4.49693
R1031 bias1.n131 bias1.t242 4.49693
R1032 bias1.n132 bias1.t309 4.49693
R1033 bias1.n132 bias1.t844 4.49693
R1034 bias1.n132 bias1.t581 4.49693
R1035 bias1.n132 bias1.t42 4.49693
R1036 bias1.n132 bias1.t623 4.49693
R1037 bias1.n132 bias1.t337 4.49693
R1038 bias1.n132 bias1.t608 4.49693
R1039 bias1.n132 bias1.t382 4.49693
R1040 bias1.n133 bias1.t448 4.49693
R1041 bias1.n133 bias1.t976 4.49693
R1042 bias1.n133 bias1.t703 4.49693
R1043 bias1.n133 bias1.t1020 4.49693
R1044 bias1.n133 bias1.t740 4.49693
R1045 bias1.n133 bias1.t483 4.49693
R1046 bias1.n133 bias1.t726 4.49693
R1047 bias1.n133 bias1.t527 4.49693
R1048 bias1.n134 bias1.t524 4.49693
R1049 bias1.n134 bias1.t1119 4.49693
R1050 bias1.n134 bias1.t835 4.49693
R1051 bias1.n134 bias1.t202 4.49693
R1052 bias1.n134 bias1.t881 4.49693
R1053 bias1.n134 bias1.t257 4.49693
R1054 bias1.n134 bias1.t864 4.49693
R1055 bias1.n134 bias1.t594 4.49693
R1056 bias1.n135 bias1.t649 4.49693
R1057 bias1.n135 bias1.t59 4.49693
R1058 bias1.n135 bias1.t632 4.49693
R1059 bias1.n135 bias1.t351 4.49693
R1060 bias1.n135 bias1.t1009 4.49693
R1061 bias1.n135 bias1.t391 4.49693
R1062 bias1.n135 bias1.t91 4.49693
R1063 bias1.n135 bias1.t375 4.49693
R1064 bias1.n136 bias1.t772 4.49693
R1065 bias1.n136 bias1.t208 4.49693
R1066 bias1.n136 bias1.t754 4.49693
R1067 bias1.n136 bias1.t496 4.49693
R1068 bias1.n136 bias1.t797 4.49693
R1069 bias1.n136 bias1.t535 4.49693
R1070 bias1.n136 bias1.t245 4.49693
R1071 bias1.n136 bias1.t521 4.49693
R1072 bias1.n137 bias1.t219 4.49693
R1073 bias1.n137 bias1.t1121 4.49693
R1074 bias1.n137 bias1.t570 4.49693
R1075 bias1.n137 bias1.t287 4.49693
R1076 bias1.n137 bias1.t816 4.49693
R1077 bias1.n137 bias1.t326 4.49693
R1078 bias1.n137 bias1.t866 4.49693
R1079 bias1.n137 bias1.t308 4.49693
R1080 bias1.n138 bias1.t1208 4.49693
R1081 bias1.n138 bias1.t62 4.49693
R1082 bias1.n138 bias1.t693 4.49693
R1083 bias1.n138 bias1.t39 4.49693
R1084 bias1.n138 bias1.t954 4.49693
R1085 bias1.n138 bias1.t471 4.49693
R1086 bias1.n138 bias1.t991 4.49693
R1087 bias1.n138 bias1.t717 4.49693
R1088 bias1.n139 bias1.t975 4.49693
R1089 bias1.n139 bias1.t142 4.49693
R1090 bias1.n139 bias1.t824 4.49693
R1091 bias1.n139 bias1.t190 4.49693
R1092 bias1.n139 bias1.t1091 4.49693
R1093 bias1.n139 bias1.t167 4.49693
R1094 bias1.n139 bias1.t1137 4.49693
R1095 bias1.n139 bias1.t855 4.49693
R1096 bias1.n2 bias1.t1118 4.49693
R1097 bias1.n2 bias1.t295 4.49693
R1098 bias1.n2 bias1.t901 4.49693
R1099 bias1.n2 bias1.t342 4.49693
R1100 bias1.n2 bias1.t30 4.49693
R1101 bias1.n2 bias1.t613 4.49693
R1102 bias1.n2 bias1.t79 4.49693
R1103 bias1.n2 bias1.t648 4.49693
R1104 bias1.n2 bias1.t58 4.49693
R1105 bias1.n2 bias1.t434 4.49693
R1106 bias1.n140 bias1.t246 4.49693
R1107 bias1.n140 bias1.t783 4.49693
R1108 bias1.n140 bias1.t220 4.49693
R1109 bias1.n141 bias1.t217 4.49693
R1110 bias1.n141 bias1.t1185 4.49693
R1111 bias1.n141 bias1.t624 4.49693
R1112 bias1.n141 bias1.t1168 4.49693
R1113 bias1.n141 bias1.t878 4.49693
R1114 bias1.n141 bias1.t1210 4.49693
R1115 bias1.n141 bias1.t923 4.49693
R1116 bias1.n141 bias1.t363 4.49693
R1117 bias1.n142 bias1.t361 4.49693
R1118 bias1.n142 bias1.t55 4.49693
R1119 bias1.n142 bias1.t404 4.49693
R1120 bias1.n142 bias1.t108 4.49693
R1121 bias1.n142 bias1.t1007 4.49693
R1122 bias1.n142 bias1.t85 4.49693
R1123 bias1.n142 bias1.t1051 4.49693
R1124 bias1.n142 bias1.t432 4.49693
R1125 bias1.n143 bias1.t510 4.49693
R1126 bias1.n143 bias1.t205 4.49693
R1127 bias1.n143 bias1.t811 4.49693
R1128 bias1.n143 bias1.t261 4.49693
R1129 bias1.n143 bias1.t793 4.49693
R1130 bias1.n143 bias1.t239 4.49693
R1131 bias1.n143 bias1.t1204 4.49693
R1132 bias1.n143 bias1.t572 4.49693
R1133 bias1.n144 bias1.t635 4.49693
R1134 bias1.n144 bias1.t1179 4.49693
R1135 bias1.n144 bias1.t894 4.49693
R1136 bias1.n144 bias1.t393 4.49693
R1137 bias1.n144 bias1.t936 4.49693
R1138 bias1.n144 bias1.t659 4.49693
R1139 bias1.n144 bias1.t916 4.49693
R1140 bias1.n144 bias1.t697 4.49693
R1141 bias1.n145 bias1.t758 4.49693
R1142 bias1.n145 bias1.t118 4.49693
R1143 bias1.n145 bias1.t1022 4.49693
R1144 bias1.n145 bias1.t161 4.49693
R1145 bias1.n145 bias1.t1067 4.49693
R1146 bias1.n145 bias1.t787 4.49693
R1147 bias1.n145 bias1.t1045 4.49693
R1148 bias1.n145 bias1.t827 4.49693
R1149 bias1.n146 bias1.t822 4.49693
R1150 bias1.n146 bias1.t274 4.49693
R1151 bias1.n146 bias1.t1171 4.49693
R1152 bias1.n146 bias1.t542 4.49693
R1153 bias1.n146 bias1.t1215 4.49693
R1154 bias1.n146 bias1.t585 4.49693
R1155 bias1.n146 bias1.t1198 4.49693
R1156 bias1.n146 bias1.t908 4.49693
R1157 bias1.n147 bias1.t958 4.49693
R1158 bias1.n147 bias1.t410 4.49693
R1159 bias1.n147 bias1.t943 4.49693
R1160 bias1.n147 bias1.t671 4.49693
R1161 bias1.n147 bias1.t150 4.49693
R1162 bias1.n147 bias1.t706 4.49693
R1163 bias1.n147 bias1.t437 4.49693
R1164 bias1.n147 bias1.t690 4.49693
R1165 bias1.n148 bias1.t1097 4.49693
R1166 bias1.n148 bias1.t548 4.49693
R1167 bias1.n148 bias1.t1079 4.49693
R1168 bias1.n148 bias1.t798 4.49693
R1169 bias1.n148 bias1.t1125 4.49693
R1170 bias1.n148 bias1.t839 4.49693
R1171 bias1.n148 bias1.t575 4.49693
R1172 bias1.n148 bias1.t819 4.49693
R1173 bias1.n149 bias1.t562 4.49693
R1174 bias1.n149 bias1.t999 4.49693
R1175 bias1.n149 bias1.t458 4.49693
R1176 bias1.n149 bias1.t152 4.49693
R1177 bias1.n149 bias1.t711 4.49693
R1178 bias1.n149 bias1.t199 4.49693
R1179 bias1.n149 bias1.t748 4.49693
R1180 bias1.n149 bias1.t178 4.49693
R1181 bias1.n150 bias1.t1083 4.49693
R1182 bias1.n150 bias1.t1145 4.49693
R1183 bias1.n150 bias1.t592 4.49693
R1184 bias1.n150 bias1.t1129 4.49693
R1185 bias1.n150 bias1.t843 4.49693
R1186 bias1.n150 bias1.t350 4.49693
R1187 bias1.n150 bias1.t889 4.49693
R1188 bias1.n150 bias1.t622 4.49693
R1189 bias1.n151 bias1.t871 4.49693
R1190 bias1.n151 bias1.t20 4.49693
R1191 bias1.n151 bias1.t714 4.49693
R1192 bias1.n151 bias1.t66 4.49693
R1193 bias1.n151 bias1.t973 4.49693
R1194 bias1.n151 bias1.t46 4.49693
R1195 bias1.n151 bias1.t1016 4.49693
R1196 bias1.n151 bias1.t738 4.49693
R1197 bias1.n2 bias1.t995 4.49693
R1198 bias1.n2 bias1.t164 4.49693
R1199 bias1.n2 bias1.t777 4.49693
R1200 bias1.n2 bias1.t213 4.49693
R1201 bias1.n2 bias1.t1115 4.49693
R1202 bias1.n2 bias1.t505 4.49693
R1203 bias1.n2 bias1.t1164 4.49693
R1204 bias1.n2 bias1.t539 4.49693
R1205 bias1.n2 bias1.t1142 4.49693
R1206 bias1.n2 bias1.t319 4.49693
R1207 bias1.t5 bias1.t0 3.48118
R1208 bias1.t6 bias1.t4 2.08438
R1209 bias1.n4 bias1.n2 1.87423
R1210 bias1.n11 bias1.n10 1.85415
R1211 bias1.n23 bias1.n22 1.69903
R1212 bias1 bias1.t207 1.61298
R1213 bias1.n2 bias1.n5 1.5757
R1214 bias1.n4 bias1.n3 1.5757
R1215 bias1.n1 bias1.n0 1.5757
R1216 bias1.n7 bias1.n6 1.57458
R1217 bias1.n1 bias1.n9 1.40929
R1218 bias1.n2 bias1.n8 1.25711
R1219 bias1.n8 bias1.n21 1.23627
R1220 bias1.n21 bias1.n20 1.23627
R1221 bias1.n20 bias1.n19 1.23627
R1222 bias1.n19 bias1.n18 1.23627
R1223 bias1.n18 bias1.n17 1.23627
R1224 bias1.n17 bias1.n16 1.23627
R1225 bias1.n16 bias1.n15 1.23627
R1226 bias1.n15 bias1.n14 1.23627
R1227 bias1.n14 bias1.n13 1.23627
R1228 bias1.n13 bias1.n12 1.23627
R1229 bias1.n12 bias1.n11 1.23627
R1230 bias1.n2 bias1.n151 1.23579
R1231 bias1.n151 bias1.n150 1.23579
R1232 bias1.n150 bias1.n149 1.23579
R1233 bias1.n149 bias1.n148 1.23579
R1234 bias1.n148 bias1.n147 1.23579
R1235 bias1.n147 bias1.n146 1.23579
R1236 bias1.n146 bias1.n145 1.23579
R1237 bias1.n145 bias1.n144 1.23579
R1238 bias1.n144 bias1.n143 1.23579
R1239 bias1.n143 bias1.n142 1.23579
R1240 bias1.n142 bias1.n141 1.23579
R1241 bias1.n141 bias1.n140 1.23579
R1242 bias1.n2 bias1.n139 1.23579
R1243 bias1.n139 bias1.n138 1.23579
R1244 bias1.n138 bias1.n137 1.23579
R1245 bias1.n137 bias1.n136 1.23579
R1246 bias1.n136 bias1.n135 1.23579
R1247 bias1.n135 bias1.n134 1.23579
R1248 bias1.n134 bias1.n133 1.23579
R1249 bias1.n133 bias1.n132 1.23579
R1250 bias1.n132 bias1.n131 1.23579
R1251 bias1.n131 bias1.n130 1.23579
R1252 bias1.n130 bias1.n129 1.23579
R1253 bias1.n129 bias1.n128 1.23579
R1254 bias1.n5 bias1.n127 1.23579
R1255 bias1.n127 bias1.n126 1.23579
R1256 bias1.n126 bias1.n125 1.23579
R1257 bias1.n125 bias1.n124 1.23579
R1258 bias1.n124 bias1.n123 1.23579
R1259 bias1.n123 bias1.n122 1.23579
R1260 bias1.n122 bias1.n121 1.23579
R1261 bias1.n121 bias1.n120 1.23579
R1262 bias1.n120 bias1.n119 1.23579
R1263 bias1.n119 bias1.n118 1.23579
R1264 bias1.n118 bias1.n117 1.23579
R1265 bias1.n117 bias1.n116 1.23579
R1266 bias1.n4 bias1.n115 1.23579
R1267 bias1.n115 bias1.n114 1.23579
R1268 bias1.n114 bias1.n113 1.23579
R1269 bias1.n113 bias1.n112 1.23579
R1270 bias1.n112 bias1.n111 1.23579
R1271 bias1.n111 bias1.n110 1.23579
R1272 bias1.n110 bias1.n109 1.23579
R1273 bias1.n109 bias1.n108 1.23579
R1274 bias1.n108 bias1.n107 1.23579
R1275 bias1.n107 bias1.n106 1.23579
R1276 bias1.n106 bias1.n105 1.23579
R1277 bias1.n105 bias1.n104 1.23579
R1278 bias1.n3 bias1.n103 1.23579
R1279 bias1.n103 bias1.n102 1.23579
R1280 bias1.n102 bias1.n101 1.23579
R1281 bias1.n101 bias1.n100 1.23579
R1282 bias1.n100 bias1.n99 1.23579
R1283 bias1.n99 bias1.n98 1.23579
R1284 bias1.n98 bias1.n97 1.23579
R1285 bias1.n97 bias1.n96 1.23579
R1286 bias1.n96 bias1.n95 1.23579
R1287 bias1.n95 bias1.n94 1.23579
R1288 bias1.n94 bias1.n93 1.23579
R1289 bias1.n93 bias1.n92 1.23579
R1290 bias1.n1 bias1.n91 1.23579
R1291 bias1.n91 bias1.n90 1.23579
R1292 bias1.n90 bias1.n89 1.23579
R1293 bias1.n89 bias1.n88 1.23579
R1294 bias1.n88 bias1.n87 1.23579
R1295 bias1.n87 bias1.n86 1.23579
R1296 bias1.n86 bias1.n85 1.23579
R1297 bias1.n85 bias1.n84 1.23579
R1298 bias1.n84 bias1.n83 1.23579
R1299 bias1.n83 bias1.n82 1.23579
R1300 bias1.n82 bias1.n81 1.23579
R1301 bias1.n81 bias1.n80 1.23579
R1302 bias1.n9 bias1.n79 1.23579
R1303 bias1.n79 bias1.n78 1.23579
R1304 bias1.n78 bias1.n77 1.23579
R1305 bias1.n77 bias1.n76 1.23579
R1306 bias1.n76 bias1.n75 1.23579
R1307 bias1.n75 bias1.n74 1.23579
R1308 bias1.n74 bias1.n73 1.23579
R1309 bias1.n73 bias1.n72 1.23579
R1310 bias1.n72 bias1.n71 1.23579
R1311 bias1.n71 bias1.n70 1.23579
R1312 bias1.n70 bias1.n69 1.23579
R1313 bias1.n69 bias1.n68 1.23579
R1314 bias1.n0 bias1.n67 1.23579
R1315 bias1.n67 bias1.n66 1.23579
R1316 bias1.n66 bias1.n65 1.23579
R1317 bias1.n65 bias1.n64 1.23579
R1318 bias1.n64 bias1.n63 1.23579
R1319 bias1.n63 bias1.n62 1.23579
R1320 bias1.n62 bias1.n61 1.23579
R1321 bias1.n61 bias1.n60 1.23579
R1322 bias1.n60 bias1.n59 1.23579
R1323 bias1.n59 bias1.n58 1.23579
R1324 bias1.n58 bias1.n57 1.23579
R1325 bias1.n57 bias1.n56 1.23579
R1326 bias1.n6 bias1.n55 1.23579
R1327 bias1.n55 bias1.n54 1.23579
R1328 bias1.n54 bias1.n53 1.23579
R1329 bias1.n53 bias1.n52 1.23579
R1330 bias1.n52 bias1.n51 1.23579
R1331 bias1.n51 bias1.n50 1.23579
R1332 bias1.n50 bias1.n49 1.23579
R1333 bias1.n49 bias1.n48 1.23579
R1334 bias1.n48 bias1.n47 1.23579
R1335 bias1.n47 bias1.n46 1.23579
R1336 bias1.n46 bias1.n45 1.23579
R1337 bias1.n45 bias1.n44 1.23579
R1338 bias1.n7 bias1.n43 1.23579
R1339 bias1.n43 bias1.n42 1.23579
R1340 bias1.n42 bias1.n41 1.23579
R1341 bias1.n41 bias1.n40 1.23579
R1342 bias1.n40 bias1.n39 1.23579
R1343 bias1.n39 bias1.n38 1.23579
R1344 bias1.n38 bias1.n37 1.23579
R1345 bias1.n37 bias1.n36 1.23579
R1346 bias1.n36 bias1.n35 1.23579
R1347 bias1.n35 bias1.n34 1.23579
R1348 bias1.n34 bias1.n33 1.23579
R1349 bias1.n33 bias1.n32 1.23579
R1350 bias1.t57 bias1.n31 1.23579
R1351 bias1.n31 bias1.n30 1.23579
R1352 bias1.n30 bias1.n29 1.23579
R1353 bias1.n29 bias1.n28 1.23579
R1354 bias1.n28 bias1.n27 1.23579
R1355 bias1.n27 bias1.n26 1.23579
R1356 bias1.n26 bias1.n25 1.23579
R1357 bias1.n25 bias1.n24 1.23579
R1358 bias1.n24 bias1.n23 1.23579
R1359 bias1.t2 bias1.t5 1.21472
R1360 bias1.t1 bias1.t2 1.21472
R1361 bias1.t3 bias1.t1 1.21472
R1362 bias1.t4 bias1.t3 1.21472
R1363 bias1 bias1.n7 1.08731
R1364 bias1.n7 bias1.n1 1.08663
R1365 bias1.n1 bias1.n4 1.08663
R1366 bias1.t231 bias1.t57 0.926969
R1367 bias1.t207 bias1.t231 0.926969
R1368 VCC.n8 VCC.n7 900
R1369 VCC.n3 VCC.n0 900
R1370 VCC.n1052 VCC.n1051 900
R1371 VCC.n1045 VCC.n1044 900
R1372 VCC.n22 VCC.t4 115.674
R1373 VCC.t17 VCC.t47 62.1823
R1374 VCC.t42 VCC.t17 62.1823
R1375 VCC.t133 VCC.t42 62.1823
R1376 VCC.t73 VCC.t133 62.1823
R1377 VCC.t97 VCC.t73 62.1823
R1378 VCC.t66 VCC.t26 62.1823
R1379 VCC.t32 VCC.t66 62.1823
R1380 VCC.t15 VCC.t32 62.1823
R1381 VCC.t58 VCC.t15 62.1823
R1382 VCC.t13 VCC.t44 45.0005
R1383 VCC.t109 VCC.t13 45.0005
R1384 VCC.t45 VCC.t109 45.0005
R1385 VCC.t60 VCC.t45 45.0005
R1386 VCC.t51 VCC.t60 45.0005
R1387 VCC.t37 VCC.t28 45.0005
R1388 VCC.t28 VCC.t22 45.0005
R1389 VCC.t22 VCC.t20 45.0005
R1390 VCC.t20 VCC.t34 45.0005
R1391 VCC.n24 VCC.t97 37.8969
R1392 VCC.n25 VCC.t58 31.1605
R1393 VCC.n25 VCC.t94 31.0223
R1394 VCC.t55 VCC.n22 29.9255
R1395 VCC.n24 VCC.t51 27.4255
R1396 VCC.t26 VCC.n24 24.286
R1397 VCC.t34 VCC.n23 22.5505
R1398 VCC.n23 VCC.t55 22.4505
R1399 VCC.n24 VCC.t37 17.5755
R1400 VCC.n18 VCC.n15 14.3291
R1401 VCC.t1040 VCC.n13 12.4255
R1402 VCC.t1039 VCC.n20 11.238
R1403 VCC.t0 VCC.t1038 10.0005
R1404 VCC.t7 VCC.t2 10.0005
R1405 VCC.t6 VCC.t1039 10.0005
R1406 VCC.n1059 VCC.t1 8.28993
R1407 VCC.n1057 VCC.t1046 7.83035
R1408 VCC.t5 VCC.t11 7.5005
R1409 VCC.t1044 VCC.t6 7.5005
R1410 VCC.n1060 VCC.t1048 7.49336
R1411 VCC.t4 VCC.t1043 6.4755
R1412 VCC.n20 VCC.t1040 6.263
R1413 VCC.t8 VCC.t9 6.0255
R1414 VCC.n1056 VCC.t12 5.71641
R1415 VCC.n1056 VCC.t3 5.71641
R1416 VCC.n1061 VCC.t1045 5.71641
R1417 VCC.n1061 VCC.t1049 5.71641
R1418 VCC.n1057 VCC.t10 5.71419
R1419 VCC.n1057 VCC.t1047 5.71419
R1420 VCC.n1059 VCC.t1037 5.71419
R1421 VCC.n124 VCC.t808 5.71419
R1422 VCC.n123 VCC.t16 5.71419
R1423 VCC.n122 VCC.t798 5.71419
R1424 VCC.n121 VCC.t393 5.71419
R1425 VCC.n120 VCC.t827 5.71419
R1426 VCC.n119 VCC.t597 5.71419
R1427 VCC.n118 VCC.t149 5.71419
R1428 VCC.n117 VCC.t629 5.71419
R1429 VCC.n116 VCC.t935 5.71419
R1430 VCC.n115 VCC.t187 5.71419
R1431 VCC.n114 VCC.t927 5.71419
R1432 VCC.n113 VCC.t725 5.71419
R1433 VCC.n112 VCC.t955 5.71419
R1434 VCC.n111 VCC.t712 5.71419
R1435 VCC.n110 VCC.t206 5.71419
R1436 VCC.n109 VCC.t750 5.71419
R1437 VCC.n108 VCC.t24 5.71419
R1438 VCC.n107 VCC.t292 5.71419
R1439 VCC.n106 VCC.t40 5.71419
R1440 VCC.n105 VCC.t498 5.71419
R1441 VCC.n104 VCC.t80 5.71419
R1442 VCC.n103 VCC.t816 5.71419
R1443 VCC.n102 VCC.t308 5.71419
R1444 VCC.n101 VCC.t807 5.71419
R1445 VCC.n100 VCC.t859 5.71419
R1446 VCC.n99 VCC.t623 5.71419
R1447 VCC.n98 VCC.t174 5.71419
R1448 VCC.n97 VCC.t609 5.71419
R1449 VCC.n96 VCC.t215 5.71419
R1450 VCC.n95 VCC.t640 5.71419
R1451 VCC.n94 VCC.t427 5.71419
R1452 VCC.n93 VCC.t933 5.71419
R1453 VCC.n92 VCC.t425 5.71419
R1454 VCC.n91 VCC.t196 5.71419
R1455 VCC.n90 VCC.t410 5.71419
R1456 VCC.n89 VCC.t186 5.71419
R1457 VCC.n88 VCC.t924 5.71419
R1458 VCC.n87 VCC.t217 5.71419
R1459 VCC.n86 VCC.t954 5.71419
R1460 VCC.n85 VCC.t433 5.71419
R1461 VCC.n84 VCC.t941 5.71419
R1462 VCC.n83 VCC.t302 5.71419
R1463 VCC.n82 VCC.t512 5.71419
R1464 VCC.n81 VCC.t288 5.71419
R1465 VCC.n80 VCC.t727 5.71419
R1466 VCC.n79 VCC.t319 5.71419
R1467 VCC.n78 VCC.t76 5.71419
R1468 VCC.n77 VCC.t529 5.71419
R1469 VCC.n76 VCC.t56 5.71419
R1470 VCC.n75 VCC.t124 5.71419
R1471 VCC.n74 VCC.t854 5.71419
R1472 VCC.n73 VCC.t398 5.71419
R1473 VCC.n72 VCC.t836 5.71419
R1474 VCC.n71 VCC.t439 5.71419
R1475 VCC.n70 VCC.t884 5.71419
R1476 VCC.n69 VCC.t638 5.71419
R1477 VCC.n68 VCC.t195 5.71419
R1478 VCC.n67 VCC.t21 5.71419
R1479 VCC.n66 VCC.t991 5.71419
R1480 VCC.n65 VCC.t230 5.71419
R1481 VCC.n64 VCC.t964 5.71419
R1482 VCC.n63 VCC.t721 5.71419
R1483 VCC.n62 VCC.t1006 5.71419
R1484 VCC.n61 VCC.t755 5.71419
R1485 VCC.n60 VCC.t250 5.71419
R1486 VCC.n59 VCC.t299 5.71419
R1487 VCC.n58 VCC.t116 5.71419
R1488 VCC.n57 VCC.t329 5.71419
R1489 VCC.n56 VCC.t88 5.71419
R1490 VCC.n55 VCC.t539 5.71419
R1491 VCC.n54 VCC.t137 5.71419
R1492 VCC.n53 VCC.t872 5.71419
R1493 VCC.n52 VCC.t353 5.71419
R1494 VCC.n51 VCC.t411 5.71419
R1495 VCC.n50 VCC.t851 5.71419
R1496 VCC.n49 VCC.t662 5.71419
R1497 VCC.n48 VCC.t219 5.71419
R1498 VCC.n47 VCC.t648 5.71419
R1499 VCC.n46 VCC.t203 5.71419
R1500 VCC.n45 VCC.t686 5.71419
R1501 VCC.n44 VCC.t468 5.71419
R1502 VCC.n43 VCC.t513 5.71419
R1503 VCC.n42 VCC.t989 5.71419
R1504 VCC.n41 VCC.t781 5.71419
R1505 VCC.n40 VCC.t1019 5.71419
R1506 VCC.n39 VCC.t765 5.71419
R1507 VCC.n38 VCC.t532 5.71419
R1508 VCC.n37 VCC.t801 5.71419
R1509 VCC.n36 VCC.t566 5.71419
R1510 VCC.n35 VCC.t564 5.71419
R1511 VCC.n34 VCC.t108 5.71419
R1512 VCC.n33 VCC.t839 5.71419
R1513 VCC.n32 VCC.t150 5.71419
R1514 VCC.n31 VCC.t887 5.71419
R1515 VCC.n30 VCC.t362 5.71419
R1516 VCC.n29 VCC.t870 5.71419
R1517 VCC.n28 VCC.t678 5.71419
R1518 VCC.n27 VCC.t674 5.71419
R1519 VCC.n125 VCC.t233 5.71419
R1520 VCC.n126 VCC.t658 5.71419
R1521 VCC.n127 VCC.t944 5.71419
R1522 VCC.n128 VCC.t490 5.71419
R1523 VCC.n129 VCC.t956 5.71419
R1524 VCC.n130 VCC.t961 5.71419
R1525 VCC.n131 VCC.t168 5.71419
R1526 VCC.n132 VCC.t616 5.71419
R1527 VCC.n133 VCC.t191 5.71419
R1528 VCC.n134 VCC.t414 5.71419
R1529 VCC.n135 VCC.t147 5.71419
R1530 VCC.n136 VCC.t376 5.71419
R1531 VCC.n137 VCC.t828 5.71419
R1532 VCC.n138 VCC.t833 5.71419
R1533 VCC.n139 VCC.t99 5.71419
R1534 VCC.n140 VCC.t787 5.71419
R1535 VCC.n141 VCC.t50 5.71419
R1536 VCC.n142 VCC.t301 5.71419
R1537 VCC.n143 VCC.t68 5.71419
R1538 VCC.n144 VCC.t275 5.71419
R1539 VCC.n145 VCC.t778 5.71419
R1540 VCC.n146 VCC.t675 5.71419
R1541 VCC.n147 VCC.t970 5.71419
R1542 VCC.n148 VCC.t465 5.71419
R1543 VCC.n149 VCC.t932 5.71419
R1544 VCC.n150 VCC.t479 5.71419
R1545 VCC.n151 VCC.t949 5.71419
R1546 VCC.n152 VCC.t160 5.71419
R1547 VCC.n153 VCC.t659 5.71419
R1548 VCC.n154 VCC.t610 5.71419
R1549 VCC.n155 VCC.t181 5.71419
R1550 VCC.n156 VCC.t400 5.71419
R1551 VCC.n157 VCC.t806 5.71419
R1552 VCC.n158 VCC.t365 5.71419
R1553 VCC.n159 VCC.t584 5.71419
R1554 VCC.n160 VCC.t382 5.71419
R1555 VCC.n161 VCC.t554 5.71419
R1556 VCC.n162 VCC.t505 5.71419
R1557 VCC.n163 VCC.t35 5.71419
R1558 VCC.n164 VCC.t291 5.71419
R1559 VCC.n165 VCC.t1008 5.71419
R1560 VCC.n166 VCC.t257 5.71419
R1561 VCC.n167 VCC.t489 5.71419
R1562 VCC.n168 VCC.t277 5.71419
R1563 VCC.n169 VCC.t455 5.71419
R1564 VCC.n170 VCC.t456 5.71419
R1565 VCC.n171 VCC.t928 5.71419
R1566 VCC.n172 VCC.t188 5.71419
R1567 VCC.n173 VCC.t689 5.71419
R1568 VCC.n174 VCC.t143 5.71419
R1569 VCC.n175 VCC.t649 5.71419
R1570 VCC.n176 VCC.t162 5.71419
R1571 VCC.n177 VCC.t389 5.71419
R1572 VCC.n178 VCC.t339 5.71419
R1573 VCC.n179 VCC.t799 5.71419
R1574 VCC.n180 VCC.t355 5.71419
R1575 VCC.n181 VCC.t576 5.71419
R1576 VCC.n182 VCC.t1017 5.71419
R1577 VCC.n183 VCC.t541 5.71419
R1578 VCC.n184 VCC.t776 5.71419
R1579 VCC.n185 VCC.t559 5.71419
R1580 VCC.n186 VCC.t239 5.71419
R1581 VCC.n187 VCC.t685 5.71419
R1582 VCC.n188 VCC.t177 5.71419
R1583 VCC.n189 VCC.t475 5.71419
R1584 VCC.n190 VCC.t207 5.71419
R1585 VCC.n191 VCC.t448 5.71419
R1586 VCC.n192 VCC.t657 5.71419
R1587 VCC.n193 VCC.t458 5.71419
R1588 VCC.n194 VCC.t673 5.71419
R1589 VCC.n195 VCC.t825 5.71419
R1590 VCC.n196 VCC.t325 5.71419
R1591 VCC.n197 VCC.t553 5.71419
R1592 VCC.n198 VCC.t107 5.71419
R1593 VCC.n199 VCC.t520 5.71419
R1594 VCC.n200 VCC.t59 5.71419
R1595 VCC.n201 VCC.t531 5.71419
R1596 VCC.n202 VCC.t762 5.71419
R1597 VCC.n203 VCC.t718 5.71419
R1598 VCC.n204 VCC.t229 5.71419
R1599 VCC.n205 VCC.t729 5.71419
R1600 VCC.n206 VCC.t987 5.71419
R1601 VCC.n207 VCC.t419 5.71419
R1602 VCC.n208 VCC.t940 5.71419
R1603 VCC.n209 VCC.t202 5.71419
R1604 VCC.n210 VCC.t953 5.71419
R1605 VCC.n211 VCC.t647 5.71419
R1606 VCC.n212 VCC.t102 5.71419
R1607 VCC.n213 VCC.t615 5.71419
R1608 VCC.n214 VCC.t850 5.71419
R1609 VCC.n215 VCC.t622 5.71419
R1610 VCC.n216 VCC.t813 5.71419
R1611 VCC.n217 VCC.t72 5.71419
R1612 VCC.n218 VCC.t826 5.71419
R1613 VCC.n219 VCC.t538 5.71419
R1614 VCC.n220 VCC.t1034 5.71419
R1615 VCC.n221 VCC.t511 5.71419
R1616 VCC.n222 VCC.t742 5.71419
R1617 VCC.n223 VCC.t298 5.71419
R1618 VCC.n224 VCC.t704 5.71419
R1619 VCC.n225 VCC.t273 5.71419
R1620 VCC.n226 VCC.t719 5.71419
R1621 VCC.n328 VCC.t745 5.71419
R1622 VCC.n327 VCC.t289 5.71419
R1623 VCC.n326 VCC.t728 5.71419
R1624 VCC.n325 VCC.t320 5.71419
R1625 VCC.n324 VCC.t761 5.71419
R1626 VCC.n323 VCC.t530 5.71419
R1627 VCC.n322 VCC.t57 5.71419
R1628 VCC.n321 VCC.t545 5.71419
R1629 VCC.n320 VCC.t853 5.71419
R1630 VCC.n319 VCC.t105 5.71419
R1631 VCC.n318 VCC.t837 5.71419
R1632 VCC.n317 VCC.t651 5.71419
R1633 VCC.n316 VCC.t885 5.71419
R1634 VCC.n315 VCC.t639 5.71419
R1635 VCC.n314 VCC.t135 5.71419
R1636 VCC.n313 VCC.t670 5.71419
R1637 VCC.n312 VCC.t988 5.71419
R1638 VCC.n311 VCC.t231 5.71419
R1639 VCC.n310 VCC.t965 5.71419
R1640 VCC.n309 VCC.t446 5.71419
R1641 VCC.n308 VCC.t1007 5.71419
R1642 VCC.n307 VCC.t756 5.71419
R1643 VCC.n306 VCC.t251 5.71419
R1644 VCC.n305 VCC.t744 5.71419
R1645 VCC.n304 VCC.t785 5.71419
R1646 VCC.n303 VCC.t556 5.71419
R1647 VCC.n302 VCC.t89 5.71419
R1648 VCC.n301 VCC.t540 5.71419
R1649 VCC.n300 VCC.t138 5.71419
R1650 VCC.n299 VCC.t571 5.71419
R1651 VCC.n298 VCC.t33 5.71419
R1652 VCC.n297 VCC.t852 5.71419
R1653 VCC.n296 VCC.t588 5.71419
R1654 VCC.n295 VCC.t370 5.71419
R1655 VCC.n294 VCC.t572 5.71419
R1656 VCC.n293 VCC.t354 5.71419
R1657 VCC.n292 VCC.t113 5.71419
R1658 VCC.n291 VCC.t387 5.71419
R1659 VCC.n290 VCC.t164 5.71419
R1660 VCC.n289 VCC.t595 5.71419
R1661 VCC.n288 VCC.t145 5.71419
R1662 VCC.n287 VCC.t488 5.71419
R1663 VCC.n286 VCC.t687 5.71419
R1664 VCC.n285 VCC.t469 5.71419
R1665 VCC.n284 VCC.t926 5.71419
R1666 VCC.n283 VCC.t501 5.71419
R1667 VCC.n282 VCC.t278 5.71419
R1668 VCC.n281 VCC.t711 5.71419
R1669 VCC.n280 VCC.t261 5.71419
R1670 VCC.n279 VCC.t23 5.71419
R1671 VCC.n278 VCC.t53 5.71419
R1672 VCC.n277 VCC.t567 5.71419
R1673 VCC.n276 VCC.t39 5.71419
R1674 VCC.n275 VCC.t601 5.71419
R1675 VCC.n274 VCC.t79 5.71419
R1676 VCC.n273 VCC.t821 5.71419
R1677 VCC.n272 VCC.t367 5.71419
R1678 VCC.n271 VCC.t364 5.71419
R1679 VCC.n270 VCC.t176 5.71419
R1680 VCC.n269 VCC.t388 5.71419
R1681 VCC.n268 VCC.t25 5.71419
R1682 VCC.n267 VCC.t916 5.71419
R1683 VCC.n266 VCC.t213 5.71419
R1684 VCC.n265 VCC.t951 5.71419
R1685 VCC.n264 VCC.t421 5.71419
R1686 VCC.n263 VCC.t478 5.71419
R1687 VCC.n262 VCC.t297 5.71419
R1688 VCC.n261 VCC.t507 5.71419
R1689 VCC.n260 VCC.t285 5.71419
R1690 VCC.n259 VCC.t723 5.71419
R1691 VCC.n258 VCC.t311 5.71419
R1692 VCC.n257 VCC.t71 5.71419
R1693 VCC.n256 VCC.t518 5.71419
R1694 VCC.n255 VCC.t574 5.71419
R1695 VCC.n254 VCC.t49 5.71419
R1696 VCC.n253 VCC.t846 5.71419
R1697 VCC.n252 VCC.t386 5.71419
R1698 VCC.n251 VCC.t830 5.71419
R1699 VCC.n250 VCC.t378 5.71419
R1700 VCC.n249 VCC.t877 5.71419
R1701 VCC.n248 VCC.t632 5.71419
R1702 VCC.n247 VCC.t693 5.71419
R1703 VCC.n246 VCC.t190 5.71419
R1704 VCC.n245 VCC.t982 5.71419
R1705 VCC.n244 VCC.t224 5.71419
R1706 VCC.n243 VCC.t959 5.71419
R1707 VCC.n242 VCC.t716 5.71419
R1708 VCC.n241 VCC.t978 5.71419
R1709 VCC.n240 VCC.t751 5.71419
R1710 VCC.n239 VCC.t748 5.71419
R1711 VCC.n238 VCC.t294 5.71419
R1712 VCC.n237 VCC.t41 5.71419
R1713 VCC.n236 VCC.t326 5.71419
R1714 VCC.n235 VCC.t82 5.71419
R1715 VCC.n234 VCC.t533 5.71419
R1716 VCC.n233 VCC.t63 5.71419
R1717 VCC.n232 VCC.t867 5.71419
R1718 VCC.n231 VCC.t861 5.71419
R1719 VCC.n230 VCC.t403 5.71419
R1720 VCC.n229 VCC.t840 5.71419
R1721 VCC.n228 VCC.t573 5.71419
R1722 VCC.n329 VCC.t139 5.71419
R1723 VCC.n330 VCC.t589 5.71419
R1724 VCC.n331 VCC.t591 5.71419
R1725 VCC.n332 VCC.t777 5.71419
R1726 VCC.n333 VCC.t283 5.71419
R1727 VCC.n334 VCC.t791 5.71419
R1728 VCC.n335 VCC.t29 5.71419
R1729 VCC.n336 VCC.t743 5.71419
R1730 VCC.n337 VCC.t1009 5.71419
R1731 VCC.n338 VCC.t491 5.71419
R1732 VCC.n339 VCC.t486 5.71419
R1733 VCC.n340 VCC.t714 5.71419
R1734 VCC.n341 VCC.t460 5.71419
R1735 VCC.n342 VCC.t677 5.71419
R1736 VCC.n343 VCC.t929 5.71419
R1737 VCC.n344 VCC.t694 5.71419
R1738 VCC.n345 VCC.t886 5.71419
R1739 VCC.n346 VCC.t440 5.71419
R1740 VCC.n347 VCC.t381 5.71419
R1741 VCC.n348 VCC.t600 5.71419
R1742 VCC.n349 VCC.t114 5.71419
R1743 VCC.n350 VCC.t565 5.71419
R1744 VCC.n351 VCC.t129 5.71419
R1745 VCC.n352 VCC.t580 5.71419
R1746 VCC.n353 VCC.t763 5.71419
R1747 VCC.n354 VCC.t321 5.71419
R1748 VCC.n355 VCC.t276 5.71419
R1749 VCC.n356 VCC.t782 5.71419
R1750 VCC.n357 VCC.t1031 5.71419
R1751 VCC.n358 VCC.t466 5.71419
R1752 VCC.n359 VCC.t1002 5.71419
R1753 VCC.n360 VCC.t252 5.71419
R1754 VCC.n361 VCC.t1013 5.71419
R1755 VCC.n362 VCC.t218 5.71419
R1756 VCC.n363 VCC.t161 5.71419
R1757 VCC.n364 VCC.t663 5.71419
R1758 VCC.n365 VCC.t911 5.71419
R1759 VCC.n366 VCC.t626 5.71419
R1760 VCC.n367 VCC.t871 5.71419
R1761 VCC.n368 VCC.t136 5.71419
R1762 VCC.n369 VCC.t889 5.71419
R1763 VCC.n370 VCC.t87 5.71419
R1764 VCC.n371 VCC.t90 5.71419
R1765 VCC.n372 VCC.t557 5.71419
R1766 VCC.n373 VCC.t788 5.71419
R1767 VCC.n374 VCC.t347 5.71419
R1768 VCC.n375 VCC.t753 5.71419
R1769 VCC.n376 VCC.t307 5.71419
R1770 VCC.n377 VCC.t768 5.71419
R1771 VCC.n378 VCC.t1022 5.71419
R1772 VCC.n379 VCC.t967 5.71419
R1773 VCC.n380 VCC.t457 5.71419
R1774 VCC.n381 VCC.t994 5.71419
R1775 VCC.n382 VCC.t243 5.71419
R1776 VCC.n383 VCC.t637 5.71419
R1777 VCC.n384 VCC.t205 5.71419
R1778 VCC.n385 VCC.t437 5.71419
R1779 VCC.n386 VCC.t225 5.71419
R1780 VCC.n387 VCC.t838 5.71419
R1781 VCC.n388 VCC.t340 5.71419
R1782 VCC.n389 VCC.t855 5.71419
R1783 VCC.n390 VCC.t126 5.71419
R1784 VCC.n391 VCC.t817 5.71419
R1785 VCC.n392 VCC.t75 5.71419
R1786 VCC.n393 VCC.t318 5.71419
R1787 VCC.n394 VCC.t92 5.71419
R1788 VCC.n395 VCC.t331 5.71419
R1789 VCC.n396 VCC.t960 5.71419
R1790 VCC.n397 VCC.t452 5.71419
R1791 VCC.n398 VCC.t666 5.71419
R1792 VCC.n399 VCC.t238 5.71419
R1793 VCC.n400 VCC.t630 5.71419
R1794 VCC.n401 VCC.t199 5.71419
R1795 VCC.n402 VCC.t646 5.71419
R1796 VCC.n403 VCC.t894 5.71419
R1797 VCC.n404 VCC.t831 5.71419
R1798 VCC.n405 VCC.t335 5.71419
R1799 VCC.n406 VCC.t848 5.71419
R1800 VCC.n407 VCC.t120 5.71419
R1801 VCC.n408 VCC.t524 5.71419
R1802 VCC.n409 VCC.t67 5.71419
R1803 VCC.n410 VCC.t309 5.71419
R1804 VCC.n411 VCC.t86 5.71419
R1805 VCC.n412 VCC.t772 5.71419
R1806 VCC.n413 VCC.t179 5.71419
R1807 VCC.n414 VCC.t735 5.71419
R1808 VCC.n415 VCC.t995 5.71419
R1809 VCC.n416 VCC.t752 5.71419
R1810 VCC.n417 VCC.t948 5.71419
R1811 VCC.n418 VCC.t210 5.71419
R1812 VCC.n419 VCC.t963 5.71419
R1813 VCC.n420 VCC.t650 5.71419
R1814 VCC.n421 VCC.t180 5.71419
R1815 VCC.n422 VCC.t620 5.71419
R1816 VCC.n423 VCC.t858 5.71419
R1817 VCC.n424 VCC.t418 5.71419
R1818 VCC.n425 VCC.t819 5.71419
R1819 VCC.n426 VCC.t383 5.71419
R1820 VCC.n427 VCC.t835 5.71419
R1821 VCC.n529 VCC.t358 5.71419
R1822 VCC.n528 VCC.t862 5.71419
R1823 VCC.n527 VCC.t344 5.71419
R1824 VCC.n526 VCC.t907 5.71419
R1825 VCC.n525 VCC.t384 5.71419
R1826 VCC.n524 VCC.t155 5.71419
R1827 VCC.n523 VCC.t635 5.71419
R1828 VCC.n522 VCC.t194 5.71419
R1829 VCC.n521 VCC.t473 5.71419
R1830 VCC.n520 VCC.t679 5.71419
R1831 VCC.n519 VCC.t461 5.71419
R1832 VCC.n518 VCC.t281 5.71419
R1833 VCC.n517 VCC.t492 5.71419
R1834 VCC.n516 VCC.t271 5.71419
R1835 VCC.n515 VCC.t700 5.71419
R1836 VCC.n514 VCC.t27 5.71419
R1837 VCC.n513 VCC.t570 5.71419
R1838 VCC.n512 VCC.t792 5.71419
R1839 VCC.n511 VCC.t562 5.71419
R1840 VCC.n510 VCC.t1030 5.71419
R1841 VCC.n509 VCC.t592 5.71419
R1842 VCC.n508 VCC.t375 5.71419
R1843 VCC.n507 VCC.t811 5.71419
R1844 VCC.n506 VCC.t356 5.71419
R1845 VCC.n505 VCC.t409 5.71419
R1846 VCC.n504 VCC.t184 5.71419
R1847 VCC.n503 VCC.t667 5.71419
R1848 VCC.n502 VCC.t166 5.71419
R1849 VCC.n501 VCC.t703 5.71419
R1850 VCC.n500 VCC.t201 5.71419
R1851 VCC.n499 VCC.t938 5.71419
R1852 VCC.n498 VCC.t471 5.71419
R1853 VCC.n497 VCC.t612 5.71419
R1854 VCC.n496 VCC.t396 5.71419
R1855 VCC.n495 VCC.t599 5.71419
R1856 VCC.n494 VCC.t377 5.71419
R1857 VCC.n493 VCC.t151 5.71419
R1858 VCC.n492 VCC.t416 5.71419
R1859 VCC.n491 VCC.t193 5.71419
R1860 VCC.n490 VCC.t618 5.71419
R1861 VCC.n489 VCC.t172 5.71419
R1862 VCC.n488 VCC.t502 5.71419
R1863 VCC.n487 VCC.t710 5.71419
R1864 VCC.n486 VCC.t487 5.71419
R1865 VCC.n485 VCC.t946 5.71419
R1866 VCC.n484 VCC.t517 5.71419
R1867 VCC.n483 VCC.t38 5.71419
R1868 VCC.n482 VCC.t731 5.71419
R1869 VCC.n481 VCC.t268 5.71419
R1870 VCC.n480 VCC.t328 5.71419
R1871 VCC.n479 VCC.t83 5.71419
R1872 VCC.n478 VCC.t586 5.71419
R1873 VCC.n477 VCC.t64 5.71419
R1874 VCC.n476 VCC.t624 5.71419
R1875 VCC.n475 VCC.t119 5.71419
R1876 VCC.n474 VCC.t786 5.71419
R1877 VCC.n473 VCC.t394 5.71419
R1878 VCC.n472 VCC.t390 5.71419
R1879 VCC.n471 VCC.t209 5.71419
R1880 VCC.n470 VCC.t428 5.71419
R1881 VCC.n469 VCC.t197 5.71419
R1882 VCC.n468 VCC.t936 5.71419
R1883 VCC.n467 VCC.t175 5.71419
R1884 VCC.n466 VCC.t975 5.71419
R1885 VCC.n465 VCC.t450 5.71419
R1886 VCC.n464 VCC.t497 5.71419
R1887 VCC.n463 VCC.t314 5.71419
R1888 VCC.n462 VCC.t526 5.71419
R1889 VCC.n461 VCC.t304 5.71419
R1890 VCC.n460 VCC.t747 5.71419
R1891 VCC.n459 VCC.t338 5.71419
R1892 VCC.n458 VCC.t103 5.71419
R1893 VCC.n457 VCC.t551 5.71419
R1894 VCC.n456 VCC.t598 5.71419
R1895 VCC.n455 VCC.t77 5.71419
R1896 VCC.n454 VCC.t881 5.71419
R1897 VCC.n453 VCC.t422 5.71419
R1898 VCC.n452 VCC.t860 5.71419
R1899 VCC.n451 VCC.t401 5.71419
R1900 VCC.n450 VCC.t905 5.71419
R1901 VCC.n449 VCC.t656 5.71419
R1902 VCC.n448 VCC.t717 5.71419
R1903 VCC.n447 VCC.t211 5.71419
R1904 VCC.n446 VCC.t979 5.71419
R1905 VCC.n445 VCC.t245 5.71419
R1906 VCC.n444 VCC.t996 5.71419
R1907 VCC.n443 VCC.t736 5.71419
R1908 VCC.n442 VCC.t1026 5.71419
R1909 VCC.n441 VCC.t774 5.71419
R1910 VCC.n440 VCC.t771 5.71419
R1911 VCC.n439 VCC.t310 5.71419
R1912 VCC.n438 VCC.t69 5.71419
R1913 VCC.n437 VCC.t349 5.71419
R1914 VCC.n436 VCC.t121 5.71419
R1915 VCC.n435 VCC.t560 5.71419
R1916 VCC.n434 VCC.t96 5.71419
R1917 VCC.n433 VCC.t897 5.71419
R1918 VCC.n432 VCC.t895 5.71419
R1919 VCC.n431 VCC.t430 5.71419
R1920 VCC.n430 VCC.t875 5.71419
R1921 VCC.n429 VCC.t496 5.71419
R1922 VCC.n530 VCC.t1032 5.71419
R1923 VCC.n531 VCC.t508 5.71419
R1924 VCC.n532 VCC.t510 5.71419
R1925 VCC.n533 VCC.t692 5.71419
R1926 VCC.n534 VCC.t198 5.71419
R1927 VCC.n535 VCC.t702 5.71419
R1928 VCC.n536 VCC.t952 5.71419
R1929 VCC.n537 VCC.t664 5.71419
R1930 VCC.n538 VCC.t917 5.71419
R1931 VCC.n539 VCC.t405 5.71419
R1932 VCC.n540 VCC.t407 5.71419
R1933 VCC.n541 VCC.t625 5.71419
R1934 VCC.n542 VCC.t372 5.71419
R1935 VCC.n543 VCC.t590 5.71419
R1936 VCC.n544 VCC.t822 5.71419
R1937 VCC.n545 VCC.t604 5.71419
R1938 VCC.n546 VCC.t790 5.71419
R1939 VCC.n547 VCC.t348 5.71419
R1940 VCC.n548 VCC.t296 5.71419
R1941 VCC.n549 VCC.t519 5.71419
R1942 VCC.n550 VCC.t976 5.71419
R1943 VCC.n551 VCC.t485 5.71419
R1944 VCC.n552 VCC.t1025 5.71419
R1945 VCC.n553 VCC.t504 5.71419
R1946 VCC.n554 VCC.t672 5.71419
R1947 VCC.n555 VCC.t244 5.71419
R1948 VCC.n556 VCC.t192 5.71419
R1949 VCC.n557 VCC.t695 5.71419
R1950 VCC.n558 VCC.t937 5.71419
R1951 VCC.n559 VCC.t380 5.71419
R1952 VCC.n560 VCC.t903 5.71419
R1953 VCC.n561 VCC.t165 5.71419
R1954 VCC.n562 VCC.t920 5.71419
R1955 VCC.n563 VCC.t111 5.71419
R1956 VCC.n564 VCC.t52 5.71419
R1957 VCC.n565 VCC.t581 5.71419
R1958 VCC.n566 VCC.t810 5.71419
R1959 VCC.n567 VCC.t542 5.71419
R1960 VCC.n568 VCC.t780 5.71419
R1961 VCC.n569 VCC.t1029 5.71419
R1962 VCC.n570 VCC.t795 5.71419
R1963 VCC.n571 VCC.t1000 5.71419
R1964 VCC.n572 VCC.t984 5.71419
R1965 VCC.n573 VCC.t482 5.71419
R1966 VCC.n574 VCC.t699 5.71419
R1967 VCC.n575 VCC.t270 5.71419
R1968 VCC.n576 VCC.t661 5.71419
R1969 VCC.n577 VCC.t236 5.71419
R1970 VCC.n578 VCC.t681 5.71419
R1971 VCC.n579 VCC.t930 5.71419
R1972 VCC.n580 VCC.t873 5.71419
R1973 VCC.n581 VCC.t369 5.71419
R1974 VCC.n582 VCC.t892 5.71419
R1975 VCC.n583 VCC.t156 5.71419
R1976 VCC.n584 VCC.t555 5.71419
R1977 VCC.n585 VCC.t118 5.71419
R1978 VCC.n586 VCC.t343 5.71419
R1979 VCC.n587 VCC.t131 5.71419
R1980 VCC.n588 VCC.t757 5.71419
R1981 VCC.n589 VCC.t263 5.71419
R1982 VCC.n590 VCC.t769 5.71419
R1983 VCC.n591 VCC.t1023 5.71419
R1984 VCC.n592 VCC.t730 5.71419
R1985 VCC.n593 VCC.t992 5.71419
R1986 VCC.n594 VCC.t241 5.71419
R1987 VCC.n595 VCC.t985 5.71419
R1988 VCC.n596 VCC.t253 5.71419
R1989 VCC.n597 VCC.t997 5.71419
R1990 VCC.n598 VCC.t474 5.71419
R1991 VCC.n599 VCC.t696 5.71419
R1992 VCC.n600 VCC.t260 5.71419
R1993 VCC.n601 VCC.t654 5.71419
R1994 VCC.n602 VCC.t228 5.71419
R1995 VCC.n603 VCC.t669 5.71419
R1996 VCC.n604 VCC.t922 5.71419
R1997 VCC.n605 VCC.t866 5.71419
R1998 VCC.n606 VCC.t359 5.71419
R1999 VCC.n607 VCC.t883 5.71419
R2000 VCC.n608 VCC.t144 5.71419
R2001 VCC.n609 VCC.t550 5.71419
R2002 VCC.n610 VCC.t98 5.71419
R2003 VCC.n611 VCC.t337 5.71419
R2004 VCC.n612 VCC.t123 5.71419
R2005 VCC.n613 VCC.t797 5.71419
R2006 VCC.n614 VCC.t256 5.71419
R2007 VCC.n615 VCC.t760 5.71419
R2008 VCC.n616 VCC.t1015 5.71419
R2009 VCC.n617 VCC.t775 5.71419
R2010 VCC.n618 VCC.t974 5.71419
R2011 VCC.n619 VCC.t237 5.71419
R2012 VCC.n620 VCC.t998 5.71419
R2013 VCC.n621 VCC.t683 5.71419
R2014 VCC.n622 VCC.t200 5.71419
R2015 VCC.n623 VCC.t644 5.71419
R2016 VCC.n624 VCC.t893 5.71419
R2017 VCC.n625 VCC.t445 5.71419
R2018 VCC.n626 VCC.t844 5.71419
R2019 VCC.n627 VCC.t406 5.71419
R2020 VCC.n628 VCC.t868 5.71419
R2021 VCC.n730 VCC.t969 5.71419
R2022 VCC.n729 VCC.t495 5.71419
R2023 VCC.n728 VCC.t945 5.71419
R2024 VCC.n727 VCC.t523 5.71419
R2025 VCC.n726 VCC.t980 5.71419
R2026 VCC.n725 VCC.t746 5.71419
R2027 VCC.n724 VCC.t290 5.71419
R2028 VCC.n723 VCC.t773 5.71419
R2029 VCC.n722 VCC.t95 5.71419
R2030 VCC.n721 VCC.t317 5.71419
R2031 VCC.n720 VCC.t74 5.71419
R2032 VCC.n719 VCC.t878 5.71419
R2033 VCC.n718 VCC.t125 5.71419
R2034 VCC.n717 VCC.t856 5.71419
R2035 VCC.n716 VCC.t341 5.71419
R2036 VCC.n715 VCC.t901 5.71419
R2037 VCC.n714 VCC.t226 5.71419
R2038 VCC.n713 VCC.t436 5.71419
R2039 VCC.n712 VCC.t204 5.71419
R2040 VCC.n711 VCC.t636 5.71419
R2041 VCC.n710 VCC.t242 5.71419
R2042 VCC.n709 VCC.t993 5.71419
R2043 VCC.n708 VCC.t454 5.71419
R2044 VCC.n707 VCC.t966 5.71419
R2045 VCC.n706 VCC.t1021 5.71419
R2046 VCC.n705 VCC.t767 5.71419
R2047 VCC.n704 VCC.t305 5.71419
R2048 VCC.n703 VCC.t754 5.71419
R2049 VCC.n702 VCC.t345 5.71419
R2050 VCC.n701 VCC.t789 5.71419
R2051 VCC.n700 VCC.t547 5.71419
R2052 VCC.n699 VCC.t91 5.71419
R2053 VCC.n698 VCC.t957 5.71419
R2054 VCC.n697 VCC.t713 5.71419
R2055 VCC.n696 VCC.t943 5.71419
R2056 VCC.n695 VCC.t698 5.71419
R2057 VCC.n694 VCC.t477 5.71419
R2058 VCC.n693 VCC.t732 5.71419
R2059 VCC.n692 VCC.t506 5.71419
R2060 VCC.n691 VCC.t968 5.71419
R2061 VCC.n690 VCC.t494 5.71419
R2062 VCC.n689 VCC.t823 5.71419
R2063 VCC.n688 VCC.t61 5.71419
R2064 VCC.n687 VCC.t805 5.71419
R2065 VCC.n686 VCC.t300 5.71419
R2066 VCC.n685 VCC.t843 5.71419
R2067 VCC.n684 VCC.t606 5.71419
R2068 VCC.n683 VCC.t93 5.71419
R2069 VCC.n682 VCC.t594 5.71419
R2070 VCC.n681 VCC.t641 5.71419
R2071 VCC.n680 VCC.t420 5.71419
R2072 VCC.n679 VCC.t934 5.71419
R2073 VCC.n678 VCC.t412 5.71419
R2074 VCC.n677 VCC.t972 5.71419
R2075 VCC.n676 VCC.t447 5.71419
R2076 VCC.n675 VCC.t221 5.71419
R2077 VCC.n674 VCC.t708 5.71419
R2078 VCC.n673 VCC.t707 5.71419
R2079 VCC.n672 VCC.t528 5.71419
R2080 VCC.n671 VCC.t740 5.71419
R2081 VCC.n670 VCC.t514 5.71419
R2082 VCC.n669 VCC.t293 5.71419
R2083 VCC.n668 VCC.t543 5.71419
R2084 VCC.n667 VCC.t323 5.71419
R2085 VCC.n666 VCC.t764 5.71419
R2086 VCC.n665 VCC.t818 5.71419
R2087 VCC.n664 VCC.t633 5.71419
R2088 VCC.n663 VCC.t857 5.71419
R2089 VCC.n662 VCC.t607 5.71419
R2090 VCC.n661 VCC.t115 5.71419
R2091 VCC.n660 VCC.t653 5.71419
R2092 VCC.n659 VCC.t442 5.71419
R2093 VCC.n658 VCC.t888 5.71419
R2094 VCC.n657 VCC.t947 5.71419
R2095 VCC.n656 VCC.t424 5.71419
R2096 VCC.n655 VCC.t246 5.71419
R2097 VCC.n654 VCC.t734 5.71419
R2098 VCC.n653 VCC.t234 5.71419
R2099 VCC.n652 VCC.t722 5.71419
R2100 VCC.n651 VCC.t264 5.71419
R2101 VCC.n650 VCC.t1011 5.71419
R2102 VCC.n649 VCC.t65 5.71419
R2103 VCC.n648 VCC.t522 5.71419
R2104 VCC.n647 VCC.t350 5.71419
R2105 VCC.n646 VCC.t558 5.71419
R2106 VCC.n645 VCC.t333 5.71419
R2107 VCC.n644 VCC.t100 5.71419
R2108 VCC.n643 VCC.t373 5.71419
R2109 VCC.n642 VCC.t141 5.71419
R2110 VCC.n641 VCC.t140 5.71419
R2111 VCC.n640 VCC.t627 5.71419
R2112 VCC.n639 VCC.t415 5.71419
R2113 VCC.n638 VCC.t665 5.71419
R2114 VCC.n637 VCC.t451 5.71419
R2115 VCC.n636 VCC.t900 5.71419
R2116 VCC.n635 VCC.t438 5.71419
R2117 VCC.n634 VCC.t258 5.71419
R2118 VCC.n633 VCC.t254 5.71419
R2119 VCC.n632 VCC.t741 5.71419
R2120 VCC.n631 VCC.t240 5.71419
R2121 VCC.n630 VCC.t417 5.71419
R2122 VCC.n731 VCC.t939 5.71419
R2123 VCC.n732 VCC.t431 5.71419
R2124 VCC.n733 VCC.t435 5.71419
R2125 VCC.n734 VCC.t603 5.71419
R2126 VCC.n735 VCC.t101 5.71419
R2127 VCC.n736 VCC.t614 5.71419
R2128 VCC.n737 VCC.t849 5.71419
R2129 VCC.n738 VCC.t583 5.71419
R2130 VCC.n739 VCC.t812 5.71419
R2131 VCC.n740 VCC.t313 5.71419
R2132 VCC.n741 VCC.t316 5.71419
R2133 VCC.n742 VCC.t537 5.71419
R2134 VCC.n743 VCC.t287 5.71419
R2135 VCC.n744 VCC.t509 5.71419
R2136 VCC.n745 VCC.t737 5.71419
R2137 VCC.n746 VCC.t521 5.71419
R2138 VCC.n747 VCC.t701 5.71419
R2139 VCC.n748 VCC.t274 5.71419
R2140 VCC.n749 VCC.t208 5.71419
R2141 VCC.n750 VCC.t444 5.71419
R2142 VCC.n751 VCC.t918 5.71419
R2143 VCC.n752 VCC.t404 5.71419
R2144 VCC.n753 VCC.t914 5.71419
R2145 VCC.n754 VCC.t423 5.71419
R2146 VCC.n755 VCC.t587 5.71419
R2147 VCC.n756 VCC.t157 5.71419
R2148 VCC.n757 VCC.t84 5.71419
R2149 VCC.n758 VCC.t608 5.71419
R2150 VCC.n759 VCC.t832 5.71419
R2151 VCC.n760 VCC.t295 5.71419
R2152 VCC.n761 VCC.t804 5.71419
R2153 VCC.n762 VCC.t54 5.71419
R2154 VCC.n763 VCC.t814 5.71419
R2155 VCC.n764 VCC.t1024 5.71419
R2156 VCC.n765 VCC.t962 5.71419
R2157 VCC.n766 VCC.t503 5.71419
R2158 VCC.n767 VCC.t726 5.71419
R2159 VCC.n768 VCC.t467 5.71419
R2160 VCC.n769 VCC.t691 5.71419
R2161 VCC.n770 VCC.t915 5.71419
R2162 VCC.n771 VCC.t705 5.71419
R2163 VCC.n772 VCC.t902 5.71419
R2164 VCC.n773 VCC.t904 5.71419
R2165 VCC.n774 VCC.t397 5.71419
R2166 VCC.n775 VCC.t613 5.71419
R2167 VCC.n776 VCC.t185 5.71419
R2168 VCC.n777 VCC.t579 5.71419
R2169 VCC.n778 VCC.t142 5.71419
R2170 VCC.n779 VCC.t593 5.71419
R2171 VCC.n780 VCC.t824 5.71419
R2172 VCC.n781 VCC.t783 5.71419
R2173 VCC.n782 VCC.t286 5.71419
R2174 VCC.n783 VCC.t796 5.71419
R2175 VCC.n784 VCC.t46 5.71419
R2176 VCC.n785 VCC.t481 5.71419
R2177 VCC.n786 VCC.t1014 5.71419
R2178 VCC.n787 VCC.t269 5.71419
R2179 VCC.n788 VCC.t1027 5.71419
R2180 VCC.n789 VCC.t544 5.71419
R2181 VCC.n790 VCC.t182 5.71419
R2182 VCC.n791 VCC.t682 5.71419
R2183 VCC.n792 VCC.t913 5.71419
R2184 VCC.n793 VCC.t643 5.71419
R2185 VCC.n794 VCC.t891 5.71419
R2186 VCC.n795 VCC.t154 5.71419
R2187 VCC.n796 VCC.t908 5.71419
R2188 VCC.n797 VCC.t169 5.71419
R2189 VCC.n798 VCC.t1016 5.71419
R2190 VCC.n799 VCC.t493 5.71419
R2191 VCC.n800 VCC.t720 5.71419
R2192 VCC.n801 VCC.t282 5.71419
R2193 VCC.n802 VCC.t684 5.71419
R2194 VCC.n803 VCC.t178 5.71419
R2195 VCC.n804 VCC.t697 5.71419
R2196 VCC.n805 VCC.t942 5.71419
R2197 VCC.n806 VCC.t896 5.71419
R2198 VCC.n807 VCC.t385 5.71419
R2199 VCC.n808 VCC.t910 5.71419
R2200 VCC.n809 VCC.t170 5.71419
R2201 VCC.n810 VCC.t569 5.71419
R2202 VCC.n811 VCC.t134 5.71419
R2203 VCC.n812 VCC.t361 5.71419
R2204 VCC.n813 VCC.t146 5.71419
R2205 VCC.n814 VCC.t815 5.71419
R2206 VCC.n815 VCC.t280 5.71419
R2207 VCC.n816 VCC.t784 5.71419
R2208 VCC.n817 VCC.t1036 5.71419
R2209 VCC.n818 VCC.t800 5.71419
R2210 VCC.n819 VCC.t1005 5.71419
R2211 VCC.n820 VCC.t259 5.71419
R2212 VCC.n821 VCC.t1018 5.71419
R2213 VCC.n822 VCC.t706 5.71419
R2214 VCC.n823 VCC.t227 5.71419
R2215 VCC.n824 VCC.t668 5.71419
R2216 VCC.n825 VCC.t921 5.71419
R2217 VCC.n826 VCC.t463 5.71419
R2218 VCC.n827 VCC.t880 5.71419
R2219 VCC.n828 VCC.t432 5.71419
R2220 VCC.n829 VCC.t898 5.71419
R2221 VCC.n931 VCC.t977 5.71419
R2222 VCC.n930 VCC.t516 5.71419
R2223 VCC.n929 VCC.t990 5.71419
R2224 VCC.n928 VCC.t549 5.71419
R2225 VCC.n927 VCC.t1020 5.71419
R2226 VCC.n926 VCC.t766 5.71419
R2227 VCC.n925 VCC.t306 5.71419
R2228 VCC.n924 VCC.t802 5.71419
R2229 VCC.n923 VCC.t130 5.71419
R2230 VCC.n922 VCC.t342 5.71419
R2231 VCC.n921 VCC.t117 5.71419
R2232 VCC.n920 VCC.t906 5.71419
R2233 VCC.n919 VCC.t152 5.71419
R2234 VCC.n918 VCC.t890 5.71419
R2235 VCC.n917 VCC.t366 5.71419
R2236 VCC.n916 VCC.t931 5.71419
R2237 VCC.n915 VCC.t248 5.71419
R2238 VCC.n914 VCC.t459 5.71419
R2239 VCC.n913 VCC.t235 5.71419
R2240 VCC.n912 VCC.t660 5.71419
R2241 VCC.n911 VCC.t265 5.71419
R2242 VCC.n910 VCC.t1012 5.71419
R2243 VCC.n909 VCC.t480 5.71419
R2244 VCC.n908 VCC.t1001 5.71419
R2245 VCC.n907 VCC.t43 5.71419
R2246 VCC.n906 VCC.t794 5.71419
R2247 VCC.n905 VCC.t334 5.71419
R2248 VCC.n904 VCC.t779 5.71419
R2249 VCC.n903 VCC.t374 5.71419
R2250 VCC.n902 VCC.t809 5.71419
R2251 VCC.n901 VCC.t578 5.71419
R2252 VCC.n900 VCC.t128 5.71419
R2253 VCC.n899 VCC.t865 5.71419
R2254 VCC.n898 VCC.t621 5.71419
R2255 VCC.n897 VCC.t842 5.71419
R2256 VCC.n896 VCC.t611 5.71419
R2257 VCC.n895 VCC.t392 5.71419
R2258 VCC.n894 VCC.t642 5.71419
R2259 VCC.n893 VCC.t429 5.71419
R2260 VCC.n892 VCC.t874 5.71419
R2261 VCC.n891 VCC.t413 5.71419
R2262 VCC.n890 VCC.t738 5.71419
R2263 VCC.n889 VCC.t971 5.71419
R2264 VCC.n888 VCC.t724 5.71419
R2265 VCC.n887 VCC.t220 5.71419
R2266 VCC.n886 VCC.t758 5.71419
R2267 VCC.n885 VCC.t527 5.71419
R2268 VCC.n884 VCC.t981 5.71419
R2269 VCC.n883 VCC.t515 5.71419
R2270 VCC.n882 VCC.t561 5.71419
R2271 VCC.n881 VCC.t336 5.71419
R2272 VCC.n880 VCC.t834 5.71419
R2273 VCC.n879 VCC.t322 5.71419
R2274 VCC.n878 VCC.t879 5.71419
R2275 VCC.n877 VCC.t357 5.71419
R2276 VCC.n876 VCC.t112 5.71419
R2277 VCC.n875 VCC.t619 5.71419
R2278 VCC.n874 VCC.t617 5.71419
R2279 VCC.n873 VCC.t453 5.71419
R2280 VCC.n872 VCC.t652 5.71419
R2281 VCC.n871 VCC.t441 5.71419
R2282 VCC.n870 VCC.t214 5.71419
R2283 VCC.n869 VCC.t472 5.71419
R2284 VCC.n868 VCC.t247 5.71419
R2285 VCC.n867 VCC.t680 5.71419
R2286 VCC.n866 VCC.t733 5.71419
R2287 VCC.n865 VCC.t552 5.71419
R2288 VCC.n864 VCC.t770 5.71419
R2289 VCC.n863 VCC.t535 5.71419
R2290 VCC.n862 VCC.t1010 5.71419
R2291 VCC.n861 VCC.t546 5.71419
R2292 VCC.n860 VCC.t351 5.71419
R2293 VCC.n859 VCC.t793 5.71419
R2294 VCC.n858 VCC.t845 5.71419
R2295 VCC.n857 VCC.t332 5.71419
R2296 VCC.n856 VCC.t158 5.71419
R2297 VCC.n855 VCC.t645 5.71419
R2298 VCC.n854 VCC.t110 5.71419
R2299 VCC.n853 VCC.t628 5.71419
R2300 VCC.n852 VCC.t183 5.71419
R2301 VCC.n851 VCC.t919 5.71419
R2302 VCC.n850 VCC.t973 5.71419
R2303 VCC.n849 VCC.t449 5.71419
R2304 VCC.n848 VCC.t272 5.71419
R2305 VCC.n847 VCC.t484 5.71419
R2306 VCC.n846 VCC.t255 5.71419
R2307 VCC.n845 VCC.t1004 5.71419
R2308 VCC.n844 VCC.t266 5.71419
R2309 VCC.n843 VCC.t1035 5.71419
R2310 VCC.n842 VCC.t1033 5.71419
R2311 VCC.n841 VCC.t548 5.71419
R2312 VCC.n840 VCC.t327 5.71419
R2313 VCC.n839 VCC.t582 5.71419
R2314 VCC.n838 VCC.t360 5.71419
R2315 VCC.n837 VCC.t803 5.71419
R2316 VCC.n836 VCC.t346 5.71419
R2317 VCC.n835 VCC.t171 5.71419
R2318 VCC.n834 VCC.t167 5.71419
R2319 VCC.n833 VCC.t655 5.71419
R2320 VCC.n832 VCC.t153 5.71419
R2321 VCC.n831 VCC.t841 5.71419
R2322 VCC.n932 VCC.t402 5.71419
R2323 VCC.n933 VCC.t864 5.71419
R2324 VCC.n934 VCC.t863 5.71419
R2325 VCC.n935 VCC.t62 5.71419
R2326 VCC.n936 VCC.t534 5.71419
R2327 VCC.n937 VCC.t81 5.71419
R2328 VCC.n938 VCC.t324 5.71419
R2329 VCC.n939 VCC.t30 5.71419
R2330 VCC.n940 VCC.t267 5.71419
R2331 VCC.n941 VCC.t749 5.71419
R2332 VCC.n942 VCC.t739 5.71419
R2333 VCC.n943 VCC.t1003 5.71419
R2334 VCC.n944 VCC.t715 5.71419
R2335 VCC.n945 VCC.t958 5.71419
R2336 VCC.n946 VCC.t223 5.71419
R2337 VCC.n947 VCC.t983 5.71419
R2338 VCC.n948 VCC.t189 5.71419
R2339 VCC.n949 VCC.t690 5.71419
R2340 VCC.n950 VCC.t631 5.71419
R2341 VCC.n951 VCC.t876 5.71419
R2342 VCC.n952 VCC.t379 5.71419
R2343 VCC.n953 VCC.t829 5.71419
R2344 VCC.n954 VCC.t395 5.71419
R2345 VCC.n955 VCC.t847 5.71419
R2346 VCC.n956 VCC.t48 5.71419
R2347 VCC.n957 VCC.t577 5.71419
R2348 VCC.n958 VCC.t525 5.71419
R2349 VCC.n959 VCC.t70 5.71419
R2350 VCC.n960 VCC.t312 5.71419
R2351 VCC.n961 VCC.t676 5.71419
R2352 VCC.n962 VCC.t284 5.71419
R2353 VCC.n963 VCC.t499 5.71419
R2354 VCC.n964 VCC.t36 5.71419
R2355 VCC.n965 VCC.t476 5.71419
R2356 VCC.n966 VCC.t426 5.71419
R2357 VCC.n967 VCC.t950 5.71419
R2358 VCC.n968 VCC.t212 5.71419
R2359 VCC.n969 VCC.t912 5.71419
R2360 VCC.n970 VCC.t173 5.71419
R2361 VCC.n971 VCC.t399 5.71419
R2362 VCC.n972 VCC.t19 5.71419
R2363 VCC.n973 VCC.t363 5.71419
R2364 VCC.n974 VCC.t368 5.71419
R2365 VCC.n975 VCC.t820 5.71419
R2366 VCC.n976 VCC.t78 5.71419
R2367 VCC.n977 VCC.t602 5.71419
R2368 VCC.n978 VCC.t14 5.71419
R2369 VCC.n979 VCC.t568 5.71419
R2370 VCC.n980 VCC.t31 5.71419
R2371 VCC.n981 VCC.t303 5.71419
R2372 VCC.n982 VCC.t262 5.71419
R2373 VCC.n983 VCC.t709 5.71419
R2374 VCC.n984 VCC.t279 5.71419
R2375 VCC.n985 VCC.t500 5.71419
R2376 VCC.n986 VCC.t925 5.71419
R2377 VCC.n987 VCC.t470 5.71419
R2378 VCC.n988 VCC.t688 5.71419
R2379 VCC.n989 VCC.t483 5.71419
R2380 VCC.n990 VCC.t148 5.71419
R2381 VCC.n991 VCC.t596 5.71419
R2382 VCC.n992 VCC.t163 5.71419
R2383 VCC.n993 VCC.t391 5.71419
R2384 VCC.n994 VCC.t127 5.71419
R2385 VCC.n995 VCC.t18 5.71419
R2386 VCC.n996 VCC.t575 5.71419
R2387 VCC.n997 VCC.t371 5.71419
R2388 VCC.n998 VCC.t585 5.71419
R2389 VCC.n999 VCC.t222 5.71419
R2390 VCC.n1000 VCC.t671 5.71419
R2391 VCC.n1001 VCC.t923 5.71419
R2392 VCC.n1002 VCC.t464 5.71419
R2393 VCC.n1003 VCC.t882 5.71419
R2394 VCC.n1004 VCC.t434 5.71419
R2395 VCC.n1005 VCC.t899 5.71419
R2396 VCC.n1006 VCC.t159 5.71419
R2397 VCC.n1007 VCC.t104 5.71419
R2398 VCC.n1008 VCC.t563 5.71419
R2399 VCC.n1009 VCC.t122 5.71419
R2400 VCC.n1010 VCC.t352 5.71419
R2401 VCC.n1011 VCC.t759 5.71419
R2402 VCC.n1012 VCC.t315 5.71419
R2403 VCC.n1013 VCC.t536 5.71419
R2404 VCC.n1014 VCC.t330 5.71419
R2405 VCC.n1015 VCC.t1028 5.71419
R2406 VCC.n1016 VCC.t462 5.71419
R2407 VCC.n1017 VCC.t999 5.71419
R2408 VCC.n1018 VCC.t249 5.71419
R2409 VCC.n1019 VCC.t986 5.71419
R2410 VCC.n1020 VCC.t216 5.71419
R2411 VCC.n1021 VCC.t443 5.71419
R2412 VCC.n1022 VCC.t232 5.71419
R2413 VCC.n1023 VCC.t909 5.71419
R2414 VCC.n1024 VCC.t408 5.71419
R2415 VCC.n1025 VCC.t869 5.71419
R2416 VCC.n1026 VCC.t132 5.71419
R2417 VCC.n1027 VCC.t634 5.71419
R2418 VCC.n1028 VCC.t85 5.71419
R2419 VCC.n1029 VCC.t605 5.71419
R2420 VCC.n1030 VCC.t106 5.71419
R2421 VCC VCC.n1063 5.09422
R2422 VCC.t1038 VCC.t1042 5.0005
R2423 VCC.t1042 VCC.t7 5.0005
R2424 VCC.n127 VCC.n126 4.63295
R2425 VCC.n229 VCC.n228 4.63295
R2426 VCC.n430 VCC.n429 4.63295
R2427 VCC.n631 VCC.n630 4.63295
R2428 VCC.n832 VCC.n831 4.63295
R2429 VCC.t1041 VCC.t0 2.5005
R2430 VCC.t2 VCC.t1044 2.5005
R2431 VCC.n629 VCC.n529 2.2255
R2432 VCC.n830 VCC.n730 2.2255
R2433 VCC.n1031 VCC.n931 2.2255
R2434 VCC.n428 VCC.n427 2.16732
R2435 VCC.n629 VCC.n628 2.16732
R2436 VCC.n830 VCC.n829 2.16732
R2437 VCC.n1031 VCC.n1030 2.16732
R2438 VCC.n227 VCC.n124 1.94545
R2439 VCC.n428 VCC.n328 1.88071
R2440 VCC.n1060 VCC.n1059 1.65712
R2441 VCC.n227 VCC.n226 1.47689
R2442 VCC.t11 VCC.t8 1.4755
R2443 VCC.t9 VCC.t1041 1.4755
R2444 VCC VCC.n1055 1.42726
R2445 VCC.t1043 VCC.t5 1.0255
R2446 VCC.n1058 VCC.n1057 0.856917
R2447 VCC.n126 VCC.n125 0.849769
R2448 VCC.n28 VCC.n27 0.849769
R2449 VCC.n29 VCC.n28 0.849769
R2450 VCC.n30 VCC.n29 0.849769
R2451 VCC.n31 VCC.n30 0.849769
R2452 VCC.n32 VCC.n31 0.849769
R2453 VCC.n33 VCC.n32 0.849769
R2454 VCC.n34 VCC.n33 0.849769
R2455 VCC.n35 VCC.n34 0.849769
R2456 VCC.n36 VCC.n35 0.849769
R2457 VCC.n37 VCC.n36 0.849769
R2458 VCC.n38 VCC.n37 0.849769
R2459 VCC.n39 VCC.n38 0.849769
R2460 VCC.n40 VCC.n39 0.849769
R2461 VCC.n41 VCC.n40 0.849769
R2462 VCC.n42 VCC.n41 0.849769
R2463 VCC.n43 VCC.n42 0.849769
R2464 VCC.n44 VCC.n43 0.849769
R2465 VCC.n45 VCC.n44 0.849769
R2466 VCC.n46 VCC.n45 0.849769
R2467 VCC.n47 VCC.n46 0.849769
R2468 VCC.n48 VCC.n47 0.849769
R2469 VCC.n49 VCC.n48 0.849769
R2470 VCC.n50 VCC.n49 0.849769
R2471 VCC.n51 VCC.n50 0.849769
R2472 VCC.n52 VCC.n51 0.849769
R2473 VCC.n53 VCC.n52 0.849769
R2474 VCC.n54 VCC.n53 0.849769
R2475 VCC.n55 VCC.n54 0.849769
R2476 VCC.n56 VCC.n55 0.849769
R2477 VCC.n57 VCC.n56 0.849769
R2478 VCC.n58 VCC.n57 0.849769
R2479 VCC.n59 VCC.n58 0.849769
R2480 VCC.n60 VCC.n59 0.849769
R2481 VCC.n61 VCC.n60 0.849769
R2482 VCC.n62 VCC.n61 0.849769
R2483 VCC.n63 VCC.n62 0.849769
R2484 VCC.n64 VCC.n63 0.849769
R2485 VCC.n65 VCC.n64 0.849769
R2486 VCC.n66 VCC.n65 0.849769
R2487 VCC.n67 VCC.n66 0.849769
R2488 VCC.n68 VCC.n67 0.849769
R2489 VCC.n69 VCC.n68 0.849769
R2490 VCC.n70 VCC.n69 0.849769
R2491 VCC.n71 VCC.n70 0.849769
R2492 VCC.n72 VCC.n71 0.849769
R2493 VCC.n73 VCC.n72 0.849769
R2494 VCC.n74 VCC.n73 0.849769
R2495 VCC.n75 VCC.n74 0.849769
R2496 VCC.n76 VCC.n75 0.849769
R2497 VCC.n77 VCC.n76 0.849769
R2498 VCC.n78 VCC.n77 0.849769
R2499 VCC.n79 VCC.n78 0.849769
R2500 VCC.n80 VCC.n79 0.849769
R2501 VCC.n81 VCC.n80 0.849769
R2502 VCC.n82 VCC.n81 0.849769
R2503 VCC.n83 VCC.n82 0.849769
R2504 VCC.n84 VCC.n83 0.849769
R2505 VCC.n85 VCC.n84 0.849769
R2506 VCC.n86 VCC.n85 0.849769
R2507 VCC.n87 VCC.n86 0.849769
R2508 VCC.n88 VCC.n87 0.849769
R2509 VCC.n89 VCC.n88 0.849769
R2510 VCC.n90 VCC.n89 0.849769
R2511 VCC.n91 VCC.n90 0.849769
R2512 VCC.n92 VCC.n91 0.849769
R2513 VCC.n93 VCC.n92 0.849769
R2514 VCC.n94 VCC.n93 0.849769
R2515 VCC.n95 VCC.n94 0.849769
R2516 VCC.n96 VCC.n95 0.849769
R2517 VCC.n97 VCC.n96 0.849769
R2518 VCC.n98 VCC.n97 0.849769
R2519 VCC.n99 VCC.n98 0.849769
R2520 VCC.n100 VCC.n99 0.849769
R2521 VCC.n101 VCC.n100 0.849769
R2522 VCC.n102 VCC.n101 0.849769
R2523 VCC.n103 VCC.n102 0.849769
R2524 VCC.n104 VCC.n103 0.849769
R2525 VCC.n105 VCC.n104 0.849769
R2526 VCC.n106 VCC.n105 0.849769
R2527 VCC.n107 VCC.n106 0.849769
R2528 VCC.n108 VCC.n107 0.849769
R2529 VCC.n109 VCC.n108 0.849769
R2530 VCC.n110 VCC.n109 0.849769
R2531 VCC.n111 VCC.n110 0.849769
R2532 VCC.n112 VCC.n111 0.849769
R2533 VCC.n113 VCC.n112 0.849769
R2534 VCC.n114 VCC.n113 0.849769
R2535 VCC.n115 VCC.n114 0.849769
R2536 VCC.n116 VCC.n115 0.849769
R2537 VCC.n117 VCC.n116 0.849769
R2538 VCC.n118 VCC.n117 0.849769
R2539 VCC.n119 VCC.n118 0.849769
R2540 VCC.n120 VCC.n119 0.849769
R2541 VCC.n121 VCC.n120 0.849769
R2542 VCC.n122 VCC.n121 0.849769
R2543 VCC.n123 VCC.n122 0.849769
R2544 VCC.n124 VCC.n123 0.849769
R2545 VCC.n427 VCC.n426 0.849769
R2546 VCC.n426 VCC.n425 0.849769
R2547 VCC.n425 VCC.n424 0.849769
R2548 VCC.n424 VCC.n423 0.849769
R2549 VCC.n423 VCC.n422 0.849769
R2550 VCC.n422 VCC.n421 0.849769
R2551 VCC.n421 VCC.n420 0.849769
R2552 VCC.n420 VCC.n419 0.849769
R2553 VCC.n419 VCC.n418 0.849769
R2554 VCC.n418 VCC.n417 0.849769
R2555 VCC.n417 VCC.n416 0.849769
R2556 VCC.n416 VCC.n415 0.849769
R2557 VCC.n415 VCC.n414 0.849769
R2558 VCC.n414 VCC.n413 0.849769
R2559 VCC.n413 VCC.n412 0.849769
R2560 VCC.n412 VCC.n411 0.849769
R2561 VCC.n411 VCC.n410 0.849769
R2562 VCC.n410 VCC.n409 0.849769
R2563 VCC.n409 VCC.n408 0.849769
R2564 VCC.n408 VCC.n407 0.849769
R2565 VCC.n407 VCC.n406 0.849769
R2566 VCC.n406 VCC.n405 0.849769
R2567 VCC.n405 VCC.n404 0.849769
R2568 VCC.n404 VCC.n403 0.849769
R2569 VCC.n403 VCC.n402 0.849769
R2570 VCC.n402 VCC.n401 0.849769
R2571 VCC.n401 VCC.n400 0.849769
R2572 VCC.n400 VCC.n399 0.849769
R2573 VCC.n399 VCC.n398 0.849769
R2574 VCC.n398 VCC.n397 0.849769
R2575 VCC.n397 VCC.n396 0.849769
R2576 VCC.n396 VCC.n395 0.849769
R2577 VCC.n395 VCC.n394 0.849769
R2578 VCC.n394 VCC.n393 0.849769
R2579 VCC.n393 VCC.n392 0.849769
R2580 VCC.n392 VCC.n391 0.849769
R2581 VCC.n391 VCC.n390 0.849769
R2582 VCC.n390 VCC.n389 0.849769
R2583 VCC.n389 VCC.n388 0.849769
R2584 VCC.n388 VCC.n387 0.849769
R2585 VCC.n387 VCC.n386 0.849769
R2586 VCC.n386 VCC.n385 0.849769
R2587 VCC.n385 VCC.n384 0.849769
R2588 VCC.n384 VCC.n383 0.849769
R2589 VCC.n383 VCC.n382 0.849769
R2590 VCC.n382 VCC.n381 0.849769
R2591 VCC.n381 VCC.n380 0.849769
R2592 VCC.n380 VCC.n379 0.849769
R2593 VCC.n379 VCC.n378 0.849769
R2594 VCC.n378 VCC.n377 0.849769
R2595 VCC.n377 VCC.n376 0.849769
R2596 VCC.n376 VCC.n375 0.849769
R2597 VCC.n375 VCC.n374 0.849769
R2598 VCC.n374 VCC.n373 0.849769
R2599 VCC.n373 VCC.n372 0.849769
R2600 VCC.n372 VCC.n371 0.849769
R2601 VCC.n371 VCC.n370 0.849769
R2602 VCC.n370 VCC.n369 0.849769
R2603 VCC.n369 VCC.n368 0.849769
R2604 VCC.n368 VCC.n367 0.849769
R2605 VCC.n367 VCC.n366 0.849769
R2606 VCC.n366 VCC.n365 0.849769
R2607 VCC.n365 VCC.n364 0.849769
R2608 VCC.n364 VCC.n363 0.849769
R2609 VCC.n363 VCC.n362 0.849769
R2610 VCC.n362 VCC.n361 0.849769
R2611 VCC.n361 VCC.n360 0.849769
R2612 VCC.n360 VCC.n359 0.849769
R2613 VCC.n359 VCC.n358 0.849769
R2614 VCC.n358 VCC.n357 0.849769
R2615 VCC.n357 VCC.n356 0.849769
R2616 VCC.n356 VCC.n355 0.849769
R2617 VCC.n355 VCC.n354 0.849769
R2618 VCC.n354 VCC.n353 0.849769
R2619 VCC.n353 VCC.n352 0.849769
R2620 VCC.n352 VCC.n351 0.849769
R2621 VCC.n351 VCC.n350 0.849769
R2622 VCC.n350 VCC.n349 0.849769
R2623 VCC.n349 VCC.n348 0.849769
R2624 VCC.n348 VCC.n347 0.849769
R2625 VCC.n347 VCC.n346 0.849769
R2626 VCC.n346 VCC.n345 0.849769
R2627 VCC.n345 VCC.n344 0.849769
R2628 VCC.n344 VCC.n343 0.849769
R2629 VCC.n343 VCC.n342 0.849769
R2630 VCC.n342 VCC.n341 0.849769
R2631 VCC.n341 VCC.n340 0.849769
R2632 VCC.n340 VCC.n339 0.849769
R2633 VCC.n339 VCC.n338 0.849769
R2634 VCC.n338 VCC.n337 0.849769
R2635 VCC.n337 VCC.n336 0.849769
R2636 VCC.n336 VCC.n335 0.849769
R2637 VCC.n335 VCC.n334 0.849769
R2638 VCC.n334 VCC.n333 0.849769
R2639 VCC.n333 VCC.n332 0.849769
R2640 VCC.n332 VCC.n331 0.849769
R2641 VCC.n331 VCC.n330 0.849769
R2642 VCC.n330 VCC.n329 0.849769
R2643 VCC.n628 VCC.n627 0.849769
R2644 VCC.n627 VCC.n626 0.849769
R2645 VCC.n626 VCC.n625 0.849769
R2646 VCC.n625 VCC.n624 0.849769
R2647 VCC.n624 VCC.n623 0.849769
R2648 VCC.n623 VCC.n622 0.849769
R2649 VCC.n622 VCC.n621 0.849769
R2650 VCC.n621 VCC.n620 0.849769
R2651 VCC.n620 VCC.n619 0.849769
R2652 VCC.n619 VCC.n618 0.849769
R2653 VCC.n618 VCC.n617 0.849769
R2654 VCC.n617 VCC.n616 0.849769
R2655 VCC.n616 VCC.n615 0.849769
R2656 VCC.n615 VCC.n614 0.849769
R2657 VCC.n614 VCC.n613 0.849769
R2658 VCC.n613 VCC.n612 0.849769
R2659 VCC.n612 VCC.n611 0.849769
R2660 VCC.n611 VCC.n610 0.849769
R2661 VCC.n610 VCC.n609 0.849769
R2662 VCC.n609 VCC.n608 0.849769
R2663 VCC.n608 VCC.n607 0.849769
R2664 VCC.n607 VCC.n606 0.849769
R2665 VCC.n606 VCC.n605 0.849769
R2666 VCC.n605 VCC.n604 0.849769
R2667 VCC.n604 VCC.n603 0.849769
R2668 VCC.n603 VCC.n602 0.849769
R2669 VCC.n602 VCC.n601 0.849769
R2670 VCC.n601 VCC.n600 0.849769
R2671 VCC.n600 VCC.n599 0.849769
R2672 VCC.n599 VCC.n598 0.849769
R2673 VCC.n598 VCC.n597 0.849769
R2674 VCC.n597 VCC.n596 0.849769
R2675 VCC.n596 VCC.n595 0.849769
R2676 VCC.n595 VCC.n594 0.849769
R2677 VCC.n594 VCC.n593 0.849769
R2678 VCC.n593 VCC.n592 0.849769
R2679 VCC.n592 VCC.n591 0.849769
R2680 VCC.n591 VCC.n590 0.849769
R2681 VCC.n590 VCC.n589 0.849769
R2682 VCC.n589 VCC.n588 0.849769
R2683 VCC.n588 VCC.n587 0.849769
R2684 VCC.n587 VCC.n586 0.849769
R2685 VCC.n586 VCC.n585 0.849769
R2686 VCC.n585 VCC.n584 0.849769
R2687 VCC.n584 VCC.n583 0.849769
R2688 VCC.n583 VCC.n582 0.849769
R2689 VCC.n582 VCC.n581 0.849769
R2690 VCC.n581 VCC.n580 0.849769
R2691 VCC.n580 VCC.n579 0.849769
R2692 VCC.n579 VCC.n578 0.849769
R2693 VCC.n578 VCC.n577 0.849769
R2694 VCC.n577 VCC.n576 0.849769
R2695 VCC.n576 VCC.n575 0.849769
R2696 VCC.n575 VCC.n574 0.849769
R2697 VCC.n574 VCC.n573 0.849769
R2698 VCC.n573 VCC.n572 0.849769
R2699 VCC.n572 VCC.n571 0.849769
R2700 VCC.n571 VCC.n570 0.849769
R2701 VCC.n570 VCC.n569 0.849769
R2702 VCC.n569 VCC.n568 0.849769
R2703 VCC.n568 VCC.n567 0.849769
R2704 VCC.n567 VCC.n566 0.849769
R2705 VCC.n566 VCC.n565 0.849769
R2706 VCC.n565 VCC.n564 0.849769
R2707 VCC.n564 VCC.n563 0.849769
R2708 VCC.n563 VCC.n562 0.849769
R2709 VCC.n562 VCC.n561 0.849769
R2710 VCC.n561 VCC.n560 0.849769
R2711 VCC.n560 VCC.n559 0.849769
R2712 VCC.n559 VCC.n558 0.849769
R2713 VCC.n558 VCC.n557 0.849769
R2714 VCC.n557 VCC.n556 0.849769
R2715 VCC.n556 VCC.n555 0.849769
R2716 VCC.n555 VCC.n554 0.849769
R2717 VCC.n554 VCC.n553 0.849769
R2718 VCC.n553 VCC.n552 0.849769
R2719 VCC.n552 VCC.n551 0.849769
R2720 VCC.n551 VCC.n550 0.849769
R2721 VCC.n550 VCC.n549 0.849769
R2722 VCC.n549 VCC.n548 0.849769
R2723 VCC.n548 VCC.n547 0.849769
R2724 VCC.n547 VCC.n546 0.849769
R2725 VCC.n546 VCC.n545 0.849769
R2726 VCC.n545 VCC.n544 0.849769
R2727 VCC.n544 VCC.n543 0.849769
R2728 VCC.n543 VCC.n542 0.849769
R2729 VCC.n542 VCC.n541 0.849769
R2730 VCC.n541 VCC.n540 0.849769
R2731 VCC.n540 VCC.n539 0.849769
R2732 VCC.n539 VCC.n538 0.849769
R2733 VCC.n538 VCC.n537 0.849769
R2734 VCC.n537 VCC.n536 0.849769
R2735 VCC.n536 VCC.n535 0.849769
R2736 VCC.n535 VCC.n534 0.849769
R2737 VCC.n534 VCC.n533 0.849769
R2738 VCC.n533 VCC.n532 0.849769
R2739 VCC.n532 VCC.n531 0.849769
R2740 VCC.n531 VCC.n530 0.849769
R2741 VCC.n829 VCC.n828 0.849769
R2742 VCC.n828 VCC.n827 0.849769
R2743 VCC.n827 VCC.n826 0.849769
R2744 VCC.n826 VCC.n825 0.849769
R2745 VCC.n825 VCC.n824 0.849769
R2746 VCC.n824 VCC.n823 0.849769
R2747 VCC.n823 VCC.n822 0.849769
R2748 VCC.n822 VCC.n821 0.849769
R2749 VCC.n821 VCC.n820 0.849769
R2750 VCC.n820 VCC.n819 0.849769
R2751 VCC.n819 VCC.n818 0.849769
R2752 VCC.n818 VCC.n817 0.849769
R2753 VCC.n817 VCC.n816 0.849769
R2754 VCC.n816 VCC.n815 0.849769
R2755 VCC.n815 VCC.n814 0.849769
R2756 VCC.n814 VCC.n813 0.849769
R2757 VCC.n813 VCC.n812 0.849769
R2758 VCC.n812 VCC.n811 0.849769
R2759 VCC.n811 VCC.n810 0.849769
R2760 VCC.n810 VCC.n809 0.849769
R2761 VCC.n809 VCC.n808 0.849769
R2762 VCC.n808 VCC.n807 0.849769
R2763 VCC.n807 VCC.n806 0.849769
R2764 VCC.n806 VCC.n805 0.849769
R2765 VCC.n805 VCC.n804 0.849769
R2766 VCC.n804 VCC.n803 0.849769
R2767 VCC.n803 VCC.n802 0.849769
R2768 VCC.n802 VCC.n801 0.849769
R2769 VCC.n801 VCC.n800 0.849769
R2770 VCC.n800 VCC.n799 0.849769
R2771 VCC.n799 VCC.n798 0.849769
R2772 VCC.n798 VCC.n797 0.849769
R2773 VCC.n797 VCC.n796 0.849769
R2774 VCC.n796 VCC.n795 0.849769
R2775 VCC.n795 VCC.n794 0.849769
R2776 VCC.n794 VCC.n793 0.849769
R2777 VCC.n793 VCC.n792 0.849769
R2778 VCC.n792 VCC.n791 0.849769
R2779 VCC.n791 VCC.n790 0.849769
R2780 VCC.n790 VCC.n789 0.849769
R2781 VCC.n789 VCC.n788 0.849769
R2782 VCC.n788 VCC.n787 0.849769
R2783 VCC.n787 VCC.n786 0.849769
R2784 VCC.n786 VCC.n785 0.849769
R2785 VCC.n785 VCC.n784 0.849769
R2786 VCC.n784 VCC.n783 0.849769
R2787 VCC.n783 VCC.n782 0.849769
R2788 VCC.n782 VCC.n781 0.849769
R2789 VCC.n781 VCC.n780 0.849769
R2790 VCC.n780 VCC.n779 0.849769
R2791 VCC.n779 VCC.n778 0.849769
R2792 VCC.n778 VCC.n777 0.849769
R2793 VCC.n777 VCC.n776 0.849769
R2794 VCC.n776 VCC.n775 0.849769
R2795 VCC.n775 VCC.n774 0.849769
R2796 VCC.n774 VCC.n773 0.849769
R2797 VCC.n773 VCC.n772 0.849769
R2798 VCC.n772 VCC.n771 0.849769
R2799 VCC.n771 VCC.n770 0.849769
R2800 VCC.n770 VCC.n769 0.849769
R2801 VCC.n769 VCC.n768 0.849769
R2802 VCC.n768 VCC.n767 0.849769
R2803 VCC.n767 VCC.n766 0.849769
R2804 VCC.n766 VCC.n765 0.849769
R2805 VCC.n765 VCC.n764 0.849769
R2806 VCC.n764 VCC.n763 0.849769
R2807 VCC.n763 VCC.n762 0.849769
R2808 VCC.n762 VCC.n761 0.849769
R2809 VCC.n761 VCC.n760 0.849769
R2810 VCC.n760 VCC.n759 0.849769
R2811 VCC.n759 VCC.n758 0.849769
R2812 VCC.n758 VCC.n757 0.849769
R2813 VCC.n757 VCC.n756 0.849769
R2814 VCC.n756 VCC.n755 0.849769
R2815 VCC.n755 VCC.n754 0.849769
R2816 VCC.n754 VCC.n753 0.849769
R2817 VCC.n753 VCC.n752 0.849769
R2818 VCC.n752 VCC.n751 0.849769
R2819 VCC.n751 VCC.n750 0.849769
R2820 VCC.n750 VCC.n749 0.849769
R2821 VCC.n749 VCC.n748 0.849769
R2822 VCC.n748 VCC.n747 0.849769
R2823 VCC.n747 VCC.n746 0.849769
R2824 VCC.n746 VCC.n745 0.849769
R2825 VCC.n745 VCC.n744 0.849769
R2826 VCC.n744 VCC.n743 0.849769
R2827 VCC.n743 VCC.n742 0.849769
R2828 VCC.n742 VCC.n741 0.849769
R2829 VCC.n741 VCC.n740 0.849769
R2830 VCC.n740 VCC.n739 0.849769
R2831 VCC.n739 VCC.n738 0.849769
R2832 VCC.n738 VCC.n737 0.849769
R2833 VCC.n737 VCC.n736 0.849769
R2834 VCC.n736 VCC.n735 0.849769
R2835 VCC.n735 VCC.n734 0.849769
R2836 VCC.n734 VCC.n733 0.849769
R2837 VCC.n733 VCC.n732 0.849769
R2838 VCC.n732 VCC.n731 0.849769
R2839 VCC.n1030 VCC.n1029 0.849769
R2840 VCC.n1029 VCC.n1028 0.849769
R2841 VCC.n1028 VCC.n1027 0.849769
R2842 VCC.n1027 VCC.n1026 0.849769
R2843 VCC.n1026 VCC.n1025 0.849769
R2844 VCC.n1025 VCC.n1024 0.849769
R2845 VCC.n1024 VCC.n1023 0.849769
R2846 VCC.n1023 VCC.n1022 0.849769
R2847 VCC.n1022 VCC.n1021 0.849769
R2848 VCC.n1021 VCC.n1020 0.849769
R2849 VCC.n1020 VCC.n1019 0.849769
R2850 VCC.n1019 VCC.n1018 0.849769
R2851 VCC.n1018 VCC.n1017 0.849769
R2852 VCC.n1017 VCC.n1016 0.849769
R2853 VCC.n1016 VCC.n1015 0.849769
R2854 VCC.n1015 VCC.n1014 0.849769
R2855 VCC.n1014 VCC.n1013 0.849769
R2856 VCC.n1013 VCC.n1012 0.849769
R2857 VCC.n1012 VCC.n1011 0.849769
R2858 VCC.n1011 VCC.n1010 0.849769
R2859 VCC.n1010 VCC.n1009 0.849769
R2860 VCC.n1009 VCC.n1008 0.849769
R2861 VCC.n1008 VCC.n1007 0.849769
R2862 VCC.n1007 VCC.n1006 0.849769
R2863 VCC.n1006 VCC.n1005 0.849769
R2864 VCC.n1005 VCC.n1004 0.849769
R2865 VCC.n1004 VCC.n1003 0.849769
R2866 VCC.n1003 VCC.n1002 0.849769
R2867 VCC.n1002 VCC.n1001 0.849769
R2868 VCC.n1001 VCC.n1000 0.849769
R2869 VCC.n1000 VCC.n999 0.849769
R2870 VCC.n999 VCC.n998 0.849769
R2871 VCC.n998 VCC.n997 0.849769
R2872 VCC.n997 VCC.n996 0.849769
R2873 VCC.n996 VCC.n995 0.849769
R2874 VCC.n995 VCC.n994 0.849769
R2875 VCC.n994 VCC.n993 0.849769
R2876 VCC.n993 VCC.n992 0.849769
R2877 VCC.n992 VCC.n991 0.849769
R2878 VCC.n991 VCC.n990 0.849769
R2879 VCC.n990 VCC.n989 0.849769
R2880 VCC.n989 VCC.n988 0.849769
R2881 VCC.n988 VCC.n987 0.849769
R2882 VCC.n987 VCC.n986 0.849769
R2883 VCC.n986 VCC.n985 0.849769
R2884 VCC.n985 VCC.n984 0.849769
R2885 VCC.n984 VCC.n983 0.849769
R2886 VCC.n983 VCC.n982 0.849769
R2887 VCC.n982 VCC.n981 0.849769
R2888 VCC.n981 VCC.n980 0.849769
R2889 VCC.n980 VCC.n979 0.849769
R2890 VCC.n979 VCC.n978 0.849769
R2891 VCC.n978 VCC.n977 0.849769
R2892 VCC.n977 VCC.n976 0.849769
R2893 VCC.n976 VCC.n975 0.849769
R2894 VCC.n975 VCC.n974 0.849769
R2895 VCC.n974 VCC.n973 0.849769
R2896 VCC.n973 VCC.n972 0.849769
R2897 VCC.n972 VCC.n971 0.849769
R2898 VCC.n971 VCC.n970 0.849769
R2899 VCC.n970 VCC.n969 0.849769
R2900 VCC.n969 VCC.n968 0.849769
R2901 VCC.n968 VCC.n967 0.849769
R2902 VCC.n967 VCC.n966 0.849769
R2903 VCC.n966 VCC.n965 0.849769
R2904 VCC.n965 VCC.n964 0.849769
R2905 VCC.n964 VCC.n963 0.849769
R2906 VCC.n963 VCC.n962 0.849769
R2907 VCC.n962 VCC.n961 0.849769
R2908 VCC.n961 VCC.n960 0.849769
R2909 VCC.n960 VCC.n959 0.849769
R2910 VCC.n959 VCC.n958 0.849769
R2911 VCC.n958 VCC.n957 0.849769
R2912 VCC.n957 VCC.n956 0.849769
R2913 VCC.n956 VCC.n955 0.849769
R2914 VCC.n955 VCC.n954 0.849769
R2915 VCC.n954 VCC.n953 0.849769
R2916 VCC.n953 VCC.n952 0.849769
R2917 VCC.n952 VCC.n951 0.849769
R2918 VCC.n951 VCC.n950 0.849769
R2919 VCC.n950 VCC.n949 0.849769
R2920 VCC.n949 VCC.n948 0.849769
R2921 VCC.n948 VCC.n947 0.849769
R2922 VCC.n947 VCC.n946 0.849769
R2923 VCC.n946 VCC.n945 0.849769
R2924 VCC.n945 VCC.n944 0.849769
R2925 VCC.n944 VCC.n943 0.849769
R2926 VCC.n943 VCC.n942 0.849769
R2927 VCC.n942 VCC.n941 0.849769
R2928 VCC.n941 VCC.n940 0.849769
R2929 VCC.n940 VCC.n939 0.849769
R2930 VCC.n939 VCC.n938 0.849769
R2931 VCC.n938 VCC.n937 0.849769
R2932 VCC.n937 VCC.n936 0.849769
R2933 VCC.n936 VCC.n935 0.849769
R2934 VCC.n935 VCC.n934 0.849769
R2935 VCC.n934 VCC.n933 0.849769
R2936 VCC.n933 VCC.n932 0.849769
R2937 VCC.n226 VCC.n225 0.789389
R2938 VCC.n225 VCC.n224 0.789389
R2939 VCC.n224 VCC.n223 0.789389
R2940 VCC.n223 VCC.n222 0.789389
R2941 VCC.n222 VCC.n221 0.789389
R2942 VCC.n221 VCC.n220 0.789389
R2943 VCC.n220 VCC.n219 0.789389
R2944 VCC.n219 VCC.n218 0.789389
R2945 VCC.n218 VCC.n217 0.789389
R2946 VCC.n217 VCC.n216 0.789389
R2947 VCC.n216 VCC.n215 0.789389
R2948 VCC.n215 VCC.n214 0.789389
R2949 VCC.n214 VCC.n213 0.789389
R2950 VCC.n213 VCC.n212 0.789389
R2951 VCC.n212 VCC.n211 0.789389
R2952 VCC.n211 VCC.n210 0.789389
R2953 VCC.n210 VCC.n209 0.789389
R2954 VCC.n209 VCC.n208 0.789389
R2955 VCC.n208 VCC.n207 0.789389
R2956 VCC.n207 VCC.n206 0.789389
R2957 VCC.n206 VCC.n205 0.789389
R2958 VCC.n205 VCC.n204 0.789389
R2959 VCC.n204 VCC.n203 0.789389
R2960 VCC.n203 VCC.n202 0.789389
R2961 VCC.n202 VCC.n201 0.789389
R2962 VCC.n201 VCC.n200 0.789389
R2963 VCC.n200 VCC.n199 0.789389
R2964 VCC.n199 VCC.n198 0.789389
R2965 VCC.n198 VCC.n197 0.789389
R2966 VCC.n197 VCC.n196 0.789389
R2967 VCC.n196 VCC.n195 0.789389
R2968 VCC.n195 VCC.n194 0.789389
R2969 VCC.n194 VCC.n193 0.789389
R2970 VCC.n193 VCC.n192 0.789389
R2971 VCC.n192 VCC.n191 0.789389
R2972 VCC.n191 VCC.n190 0.789389
R2973 VCC.n190 VCC.n189 0.789389
R2974 VCC.n189 VCC.n188 0.789389
R2975 VCC.n188 VCC.n187 0.789389
R2976 VCC.n187 VCC.n186 0.789389
R2977 VCC.n186 VCC.n185 0.789389
R2978 VCC.n185 VCC.n184 0.789389
R2979 VCC.n184 VCC.n183 0.789389
R2980 VCC.n183 VCC.n182 0.789389
R2981 VCC.n182 VCC.n181 0.789389
R2982 VCC.n181 VCC.n180 0.789389
R2983 VCC.n180 VCC.n179 0.789389
R2984 VCC.n179 VCC.n178 0.789389
R2985 VCC.n178 VCC.n177 0.789389
R2986 VCC.n177 VCC.n176 0.789389
R2987 VCC.n176 VCC.n175 0.789389
R2988 VCC.n175 VCC.n174 0.789389
R2989 VCC.n174 VCC.n173 0.789389
R2990 VCC.n173 VCC.n172 0.789389
R2991 VCC.n172 VCC.n171 0.789389
R2992 VCC.n171 VCC.n170 0.789389
R2993 VCC.n170 VCC.n169 0.789389
R2994 VCC.n169 VCC.n168 0.789389
R2995 VCC.n168 VCC.n167 0.789389
R2996 VCC.n167 VCC.n166 0.789389
R2997 VCC.n166 VCC.n165 0.789389
R2998 VCC.n165 VCC.n164 0.789389
R2999 VCC.n164 VCC.n163 0.789389
R3000 VCC.n163 VCC.n162 0.789389
R3001 VCC.n162 VCC.n161 0.789389
R3002 VCC.n161 VCC.n160 0.789389
R3003 VCC.n160 VCC.n159 0.789389
R3004 VCC.n159 VCC.n158 0.789389
R3005 VCC.n158 VCC.n157 0.789389
R3006 VCC.n157 VCC.n156 0.789389
R3007 VCC.n156 VCC.n155 0.789389
R3008 VCC.n155 VCC.n154 0.789389
R3009 VCC.n154 VCC.n153 0.789389
R3010 VCC.n153 VCC.n152 0.789389
R3011 VCC.n152 VCC.n151 0.789389
R3012 VCC.n151 VCC.n150 0.789389
R3013 VCC.n150 VCC.n149 0.789389
R3014 VCC.n149 VCC.n148 0.789389
R3015 VCC.n148 VCC.n147 0.789389
R3016 VCC.n147 VCC.n146 0.789389
R3017 VCC.n146 VCC.n145 0.789389
R3018 VCC.n145 VCC.n144 0.789389
R3019 VCC.n144 VCC.n143 0.789389
R3020 VCC.n143 VCC.n142 0.789389
R3021 VCC.n142 VCC.n141 0.789389
R3022 VCC.n141 VCC.n140 0.789389
R3023 VCC.n140 VCC.n139 0.789389
R3024 VCC.n139 VCC.n138 0.789389
R3025 VCC.n138 VCC.n137 0.789389
R3026 VCC.n137 VCC.n136 0.789389
R3027 VCC.n136 VCC.n135 0.789389
R3028 VCC.n135 VCC.n134 0.789389
R3029 VCC.n134 VCC.n133 0.789389
R3030 VCC.n133 VCC.n132 0.789389
R3031 VCC.n132 VCC.n131 0.789389
R3032 VCC.n131 VCC.n130 0.789389
R3033 VCC.n130 VCC.n129 0.789389
R3034 VCC.n129 VCC.n128 0.789389
R3035 VCC.n128 VCC.n127 0.789389
R3036 VCC.n230 VCC.n229 0.789389
R3037 VCC.n231 VCC.n230 0.789389
R3038 VCC.n232 VCC.n231 0.789389
R3039 VCC.n233 VCC.n232 0.789389
R3040 VCC.n234 VCC.n233 0.789389
R3041 VCC.n235 VCC.n234 0.789389
R3042 VCC.n236 VCC.n235 0.789389
R3043 VCC.n237 VCC.n236 0.789389
R3044 VCC.n238 VCC.n237 0.789389
R3045 VCC.n239 VCC.n238 0.789389
R3046 VCC.n240 VCC.n239 0.789389
R3047 VCC.n241 VCC.n240 0.789389
R3048 VCC.n242 VCC.n241 0.789389
R3049 VCC.n243 VCC.n242 0.789389
R3050 VCC.n244 VCC.n243 0.789389
R3051 VCC.n245 VCC.n244 0.789389
R3052 VCC.n246 VCC.n245 0.789389
R3053 VCC.n247 VCC.n246 0.789389
R3054 VCC.n248 VCC.n247 0.789389
R3055 VCC.n249 VCC.n248 0.789389
R3056 VCC.n250 VCC.n249 0.789389
R3057 VCC.n251 VCC.n250 0.789389
R3058 VCC.n252 VCC.n251 0.789389
R3059 VCC.n253 VCC.n252 0.789389
R3060 VCC.n254 VCC.n253 0.789389
R3061 VCC.n255 VCC.n254 0.789389
R3062 VCC.n256 VCC.n255 0.789389
R3063 VCC.n257 VCC.n256 0.789389
R3064 VCC.n258 VCC.n257 0.789389
R3065 VCC.n259 VCC.n258 0.789389
R3066 VCC.n260 VCC.n259 0.789389
R3067 VCC.n261 VCC.n260 0.789389
R3068 VCC.n262 VCC.n261 0.789389
R3069 VCC.n263 VCC.n262 0.789389
R3070 VCC.n264 VCC.n263 0.789389
R3071 VCC.n265 VCC.n264 0.789389
R3072 VCC.n266 VCC.n265 0.789389
R3073 VCC.n267 VCC.n266 0.789389
R3074 VCC.n268 VCC.n267 0.789389
R3075 VCC.n269 VCC.n268 0.789389
R3076 VCC.n270 VCC.n269 0.789389
R3077 VCC.n271 VCC.n270 0.789389
R3078 VCC.n272 VCC.n271 0.789389
R3079 VCC.n273 VCC.n272 0.789389
R3080 VCC.n274 VCC.n273 0.789389
R3081 VCC.n275 VCC.n274 0.789389
R3082 VCC.n276 VCC.n275 0.789389
R3083 VCC.n277 VCC.n276 0.789389
R3084 VCC.n278 VCC.n277 0.789389
R3085 VCC.n279 VCC.n278 0.789389
R3086 VCC.n280 VCC.n279 0.789389
R3087 VCC.n281 VCC.n280 0.789389
R3088 VCC.n282 VCC.n281 0.789389
R3089 VCC.n283 VCC.n282 0.789389
R3090 VCC.n284 VCC.n283 0.789389
R3091 VCC.n285 VCC.n284 0.789389
R3092 VCC.n286 VCC.n285 0.789389
R3093 VCC.n287 VCC.n286 0.789389
R3094 VCC.n288 VCC.n287 0.789389
R3095 VCC.n289 VCC.n288 0.789389
R3096 VCC.n290 VCC.n289 0.789389
R3097 VCC.n291 VCC.n290 0.789389
R3098 VCC.n292 VCC.n291 0.789389
R3099 VCC.n293 VCC.n292 0.789389
R3100 VCC.n294 VCC.n293 0.789389
R3101 VCC.n295 VCC.n294 0.789389
R3102 VCC.n296 VCC.n295 0.789389
R3103 VCC.n297 VCC.n296 0.789389
R3104 VCC.n298 VCC.n297 0.789389
R3105 VCC.n299 VCC.n298 0.789389
R3106 VCC.n300 VCC.n299 0.789389
R3107 VCC.n301 VCC.n300 0.789389
R3108 VCC.n302 VCC.n301 0.789389
R3109 VCC.n303 VCC.n302 0.789389
R3110 VCC.n304 VCC.n303 0.789389
R3111 VCC.n305 VCC.n304 0.789389
R3112 VCC.n306 VCC.n305 0.789389
R3113 VCC.n307 VCC.n306 0.789389
R3114 VCC.n308 VCC.n307 0.789389
R3115 VCC.n309 VCC.n308 0.789389
R3116 VCC.n310 VCC.n309 0.789389
R3117 VCC.n311 VCC.n310 0.789389
R3118 VCC.n312 VCC.n311 0.789389
R3119 VCC.n313 VCC.n312 0.789389
R3120 VCC.n314 VCC.n313 0.789389
R3121 VCC.n315 VCC.n314 0.789389
R3122 VCC.n316 VCC.n315 0.789389
R3123 VCC.n317 VCC.n316 0.789389
R3124 VCC.n318 VCC.n317 0.789389
R3125 VCC.n319 VCC.n318 0.789389
R3126 VCC.n320 VCC.n319 0.789389
R3127 VCC.n321 VCC.n320 0.789389
R3128 VCC.n322 VCC.n321 0.789389
R3129 VCC.n323 VCC.n322 0.789389
R3130 VCC.n324 VCC.n323 0.789389
R3131 VCC.n325 VCC.n324 0.789389
R3132 VCC.n326 VCC.n325 0.789389
R3133 VCC.n327 VCC.n326 0.789389
R3134 VCC.n328 VCC.n327 0.789389
R3135 VCC.n431 VCC.n430 0.789389
R3136 VCC.n432 VCC.n431 0.789389
R3137 VCC.n433 VCC.n432 0.789389
R3138 VCC.n434 VCC.n433 0.789389
R3139 VCC.n435 VCC.n434 0.789389
R3140 VCC.n436 VCC.n435 0.789389
R3141 VCC.n437 VCC.n436 0.789389
R3142 VCC.n438 VCC.n437 0.789389
R3143 VCC.n439 VCC.n438 0.789389
R3144 VCC.n440 VCC.n439 0.789389
R3145 VCC.n441 VCC.n440 0.789389
R3146 VCC.n442 VCC.n441 0.789389
R3147 VCC.n443 VCC.n442 0.789389
R3148 VCC.n444 VCC.n443 0.789389
R3149 VCC.n445 VCC.n444 0.789389
R3150 VCC.n446 VCC.n445 0.789389
R3151 VCC.n447 VCC.n446 0.789389
R3152 VCC.n448 VCC.n447 0.789389
R3153 VCC.n449 VCC.n448 0.789389
R3154 VCC.n450 VCC.n449 0.789389
R3155 VCC.n451 VCC.n450 0.789389
R3156 VCC.n452 VCC.n451 0.789389
R3157 VCC.n453 VCC.n452 0.789389
R3158 VCC.n454 VCC.n453 0.789389
R3159 VCC.n455 VCC.n454 0.789389
R3160 VCC.n456 VCC.n455 0.789389
R3161 VCC.n457 VCC.n456 0.789389
R3162 VCC.n458 VCC.n457 0.789389
R3163 VCC.n459 VCC.n458 0.789389
R3164 VCC.n460 VCC.n459 0.789389
R3165 VCC.n461 VCC.n460 0.789389
R3166 VCC.n462 VCC.n461 0.789389
R3167 VCC.n463 VCC.n462 0.789389
R3168 VCC.n464 VCC.n463 0.789389
R3169 VCC.n465 VCC.n464 0.789389
R3170 VCC.n466 VCC.n465 0.789389
R3171 VCC.n467 VCC.n466 0.789389
R3172 VCC.n468 VCC.n467 0.789389
R3173 VCC.n469 VCC.n468 0.789389
R3174 VCC.n470 VCC.n469 0.789389
R3175 VCC.n471 VCC.n470 0.789389
R3176 VCC.n472 VCC.n471 0.789389
R3177 VCC.n473 VCC.n472 0.789389
R3178 VCC.n474 VCC.n473 0.789389
R3179 VCC.n475 VCC.n474 0.789389
R3180 VCC.n476 VCC.n475 0.789389
R3181 VCC.n477 VCC.n476 0.789389
R3182 VCC.n478 VCC.n477 0.789389
R3183 VCC.n479 VCC.n478 0.789389
R3184 VCC.n480 VCC.n479 0.789389
R3185 VCC.n481 VCC.n480 0.789389
R3186 VCC.n482 VCC.n481 0.789389
R3187 VCC.n483 VCC.n482 0.789389
R3188 VCC.n484 VCC.n483 0.789389
R3189 VCC.n485 VCC.n484 0.789389
R3190 VCC.n486 VCC.n485 0.789389
R3191 VCC.n487 VCC.n486 0.789389
R3192 VCC.n488 VCC.n487 0.789389
R3193 VCC.n489 VCC.n488 0.789389
R3194 VCC.n490 VCC.n489 0.789389
R3195 VCC.n491 VCC.n490 0.789389
R3196 VCC.n492 VCC.n491 0.789389
R3197 VCC.n493 VCC.n492 0.789389
R3198 VCC.n494 VCC.n493 0.789389
R3199 VCC.n495 VCC.n494 0.789389
R3200 VCC.n496 VCC.n495 0.789389
R3201 VCC.n497 VCC.n496 0.789389
R3202 VCC.n498 VCC.n497 0.789389
R3203 VCC.n499 VCC.n498 0.789389
R3204 VCC.n500 VCC.n499 0.789389
R3205 VCC.n501 VCC.n500 0.789389
R3206 VCC.n502 VCC.n501 0.789389
R3207 VCC.n503 VCC.n502 0.789389
R3208 VCC.n504 VCC.n503 0.789389
R3209 VCC.n505 VCC.n504 0.789389
R3210 VCC.n506 VCC.n505 0.789389
R3211 VCC.n507 VCC.n506 0.789389
R3212 VCC.n508 VCC.n507 0.789389
R3213 VCC.n509 VCC.n508 0.789389
R3214 VCC.n510 VCC.n509 0.789389
R3215 VCC.n511 VCC.n510 0.789389
R3216 VCC.n512 VCC.n511 0.789389
R3217 VCC.n513 VCC.n512 0.789389
R3218 VCC.n514 VCC.n513 0.789389
R3219 VCC.n515 VCC.n514 0.789389
R3220 VCC.n516 VCC.n515 0.789389
R3221 VCC.n517 VCC.n516 0.789389
R3222 VCC.n518 VCC.n517 0.789389
R3223 VCC.n519 VCC.n518 0.789389
R3224 VCC.n520 VCC.n519 0.789389
R3225 VCC.n521 VCC.n520 0.789389
R3226 VCC.n522 VCC.n521 0.789389
R3227 VCC.n523 VCC.n522 0.789389
R3228 VCC.n524 VCC.n523 0.789389
R3229 VCC.n525 VCC.n524 0.789389
R3230 VCC.n526 VCC.n525 0.789389
R3231 VCC.n527 VCC.n526 0.789389
R3232 VCC.n528 VCC.n527 0.789389
R3233 VCC.n529 VCC.n528 0.789389
R3234 VCC.n632 VCC.n631 0.789389
R3235 VCC.n633 VCC.n632 0.789389
R3236 VCC.n634 VCC.n633 0.789389
R3237 VCC.n635 VCC.n634 0.789389
R3238 VCC.n636 VCC.n635 0.789389
R3239 VCC.n637 VCC.n636 0.789389
R3240 VCC.n638 VCC.n637 0.789389
R3241 VCC.n639 VCC.n638 0.789389
R3242 VCC.n640 VCC.n639 0.789389
R3243 VCC.n641 VCC.n640 0.789389
R3244 VCC.n642 VCC.n641 0.789389
R3245 VCC.n643 VCC.n642 0.789389
R3246 VCC.n644 VCC.n643 0.789389
R3247 VCC.n645 VCC.n644 0.789389
R3248 VCC.n646 VCC.n645 0.789389
R3249 VCC.n647 VCC.n646 0.789389
R3250 VCC.n648 VCC.n647 0.789389
R3251 VCC.n649 VCC.n648 0.789389
R3252 VCC.n650 VCC.n649 0.789389
R3253 VCC.n651 VCC.n650 0.789389
R3254 VCC.n652 VCC.n651 0.789389
R3255 VCC.n653 VCC.n652 0.789389
R3256 VCC.n654 VCC.n653 0.789389
R3257 VCC.n655 VCC.n654 0.789389
R3258 VCC.n656 VCC.n655 0.789389
R3259 VCC.n657 VCC.n656 0.789389
R3260 VCC.n658 VCC.n657 0.789389
R3261 VCC.n659 VCC.n658 0.789389
R3262 VCC.n660 VCC.n659 0.789389
R3263 VCC.n661 VCC.n660 0.789389
R3264 VCC.n662 VCC.n661 0.789389
R3265 VCC.n663 VCC.n662 0.789389
R3266 VCC.n664 VCC.n663 0.789389
R3267 VCC.n665 VCC.n664 0.789389
R3268 VCC.n666 VCC.n665 0.789389
R3269 VCC.n667 VCC.n666 0.789389
R3270 VCC.n668 VCC.n667 0.789389
R3271 VCC.n669 VCC.n668 0.789389
R3272 VCC.n670 VCC.n669 0.789389
R3273 VCC.n671 VCC.n670 0.789389
R3274 VCC.n672 VCC.n671 0.789389
R3275 VCC.n673 VCC.n672 0.789389
R3276 VCC.n674 VCC.n673 0.789389
R3277 VCC.n675 VCC.n674 0.789389
R3278 VCC.n676 VCC.n675 0.789389
R3279 VCC.n677 VCC.n676 0.789389
R3280 VCC.n678 VCC.n677 0.789389
R3281 VCC.n679 VCC.n678 0.789389
R3282 VCC.n680 VCC.n679 0.789389
R3283 VCC.n681 VCC.n680 0.789389
R3284 VCC.n682 VCC.n681 0.789389
R3285 VCC.n683 VCC.n682 0.789389
R3286 VCC.n684 VCC.n683 0.789389
R3287 VCC.n685 VCC.n684 0.789389
R3288 VCC.n686 VCC.n685 0.789389
R3289 VCC.n687 VCC.n686 0.789389
R3290 VCC.n688 VCC.n687 0.789389
R3291 VCC.n689 VCC.n688 0.789389
R3292 VCC.n690 VCC.n689 0.789389
R3293 VCC.n691 VCC.n690 0.789389
R3294 VCC.n692 VCC.n691 0.789389
R3295 VCC.n693 VCC.n692 0.789389
R3296 VCC.n694 VCC.n693 0.789389
R3297 VCC.n695 VCC.n694 0.789389
R3298 VCC.n696 VCC.n695 0.789389
R3299 VCC.n697 VCC.n696 0.789389
R3300 VCC.n698 VCC.n697 0.789389
R3301 VCC.n699 VCC.n698 0.789389
R3302 VCC.n700 VCC.n699 0.789389
R3303 VCC.n701 VCC.n700 0.789389
R3304 VCC.n702 VCC.n701 0.789389
R3305 VCC.n703 VCC.n702 0.789389
R3306 VCC.n704 VCC.n703 0.789389
R3307 VCC.n705 VCC.n704 0.789389
R3308 VCC.n706 VCC.n705 0.789389
R3309 VCC.n707 VCC.n706 0.789389
R3310 VCC.n708 VCC.n707 0.789389
R3311 VCC.n709 VCC.n708 0.789389
R3312 VCC.n710 VCC.n709 0.789389
R3313 VCC.n711 VCC.n710 0.789389
R3314 VCC.n712 VCC.n711 0.789389
R3315 VCC.n713 VCC.n712 0.789389
R3316 VCC.n714 VCC.n713 0.789389
R3317 VCC.n715 VCC.n714 0.789389
R3318 VCC.n716 VCC.n715 0.789389
R3319 VCC.n717 VCC.n716 0.789389
R3320 VCC.n718 VCC.n717 0.789389
R3321 VCC.n719 VCC.n718 0.789389
R3322 VCC.n720 VCC.n719 0.789389
R3323 VCC.n721 VCC.n720 0.789389
R3324 VCC.n722 VCC.n721 0.789389
R3325 VCC.n723 VCC.n722 0.789389
R3326 VCC.n724 VCC.n723 0.789389
R3327 VCC.n725 VCC.n724 0.789389
R3328 VCC.n726 VCC.n725 0.789389
R3329 VCC.n727 VCC.n726 0.789389
R3330 VCC.n728 VCC.n727 0.789389
R3331 VCC.n729 VCC.n728 0.789389
R3332 VCC.n730 VCC.n729 0.789389
R3333 VCC.n833 VCC.n832 0.789389
R3334 VCC.n834 VCC.n833 0.789389
R3335 VCC.n835 VCC.n834 0.789389
R3336 VCC.n836 VCC.n835 0.789389
R3337 VCC.n837 VCC.n836 0.789389
R3338 VCC.n838 VCC.n837 0.789389
R3339 VCC.n839 VCC.n838 0.789389
R3340 VCC.n840 VCC.n839 0.789389
R3341 VCC.n841 VCC.n840 0.789389
R3342 VCC.n842 VCC.n841 0.789389
R3343 VCC.n843 VCC.n842 0.789389
R3344 VCC.n844 VCC.n843 0.789389
R3345 VCC.n845 VCC.n844 0.789389
R3346 VCC.n846 VCC.n845 0.789389
R3347 VCC.n847 VCC.n846 0.789389
R3348 VCC.n848 VCC.n847 0.789389
R3349 VCC.n849 VCC.n848 0.789389
R3350 VCC.n850 VCC.n849 0.789389
R3351 VCC.n851 VCC.n850 0.789389
R3352 VCC.n852 VCC.n851 0.789389
R3353 VCC.n853 VCC.n852 0.789389
R3354 VCC.n854 VCC.n853 0.789389
R3355 VCC.n855 VCC.n854 0.789389
R3356 VCC.n856 VCC.n855 0.789389
R3357 VCC.n857 VCC.n856 0.789389
R3358 VCC.n858 VCC.n857 0.789389
R3359 VCC.n859 VCC.n858 0.789389
R3360 VCC.n860 VCC.n859 0.789389
R3361 VCC.n861 VCC.n860 0.789389
R3362 VCC.n862 VCC.n861 0.789389
R3363 VCC.n863 VCC.n862 0.789389
R3364 VCC.n864 VCC.n863 0.789389
R3365 VCC.n865 VCC.n864 0.789389
R3366 VCC.n866 VCC.n865 0.789389
R3367 VCC.n867 VCC.n866 0.789389
R3368 VCC.n868 VCC.n867 0.789389
R3369 VCC.n869 VCC.n868 0.789389
R3370 VCC.n870 VCC.n869 0.789389
R3371 VCC.n871 VCC.n870 0.789389
R3372 VCC.n872 VCC.n871 0.789389
R3373 VCC.n873 VCC.n872 0.789389
R3374 VCC.n874 VCC.n873 0.789389
R3375 VCC.n875 VCC.n874 0.789389
R3376 VCC.n876 VCC.n875 0.789389
R3377 VCC.n877 VCC.n876 0.789389
R3378 VCC.n878 VCC.n877 0.789389
R3379 VCC.n879 VCC.n878 0.789389
R3380 VCC.n880 VCC.n879 0.789389
R3381 VCC.n881 VCC.n880 0.789389
R3382 VCC.n882 VCC.n881 0.789389
R3383 VCC.n883 VCC.n882 0.789389
R3384 VCC.n884 VCC.n883 0.789389
R3385 VCC.n885 VCC.n884 0.789389
R3386 VCC.n886 VCC.n885 0.789389
R3387 VCC.n887 VCC.n886 0.789389
R3388 VCC.n888 VCC.n887 0.789389
R3389 VCC.n889 VCC.n888 0.789389
R3390 VCC.n890 VCC.n889 0.789389
R3391 VCC.n891 VCC.n890 0.789389
R3392 VCC.n892 VCC.n891 0.789389
R3393 VCC.n893 VCC.n892 0.789389
R3394 VCC.n894 VCC.n893 0.789389
R3395 VCC.n895 VCC.n894 0.789389
R3396 VCC.n896 VCC.n895 0.789389
R3397 VCC.n897 VCC.n896 0.789389
R3398 VCC.n898 VCC.n897 0.789389
R3399 VCC.n899 VCC.n898 0.789389
R3400 VCC.n900 VCC.n899 0.789389
R3401 VCC.n901 VCC.n900 0.789389
R3402 VCC.n902 VCC.n901 0.789389
R3403 VCC.n903 VCC.n902 0.789389
R3404 VCC.n904 VCC.n903 0.789389
R3405 VCC.n905 VCC.n904 0.789389
R3406 VCC.n906 VCC.n905 0.789389
R3407 VCC.n907 VCC.n906 0.789389
R3408 VCC.n908 VCC.n907 0.789389
R3409 VCC.n909 VCC.n908 0.789389
R3410 VCC.n910 VCC.n909 0.789389
R3411 VCC.n911 VCC.n910 0.789389
R3412 VCC.n912 VCC.n911 0.789389
R3413 VCC.n913 VCC.n912 0.789389
R3414 VCC.n914 VCC.n913 0.789389
R3415 VCC.n915 VCC.n914 0.789389
R3416 VCC.n916 VCC.n915 0.789389
R3417 VCC.n917 VCC.n916 0.789389
R3418 VCC.n918 VCC.n917 0.789389
R3419 VCC.n919 VCC.n918 0.789389
R3420 VCC.n920 VCC.n919 0.789389
R3421 VCC.n921 VCC.n920 0.789389
R3422 VCC.n922 VCC.n921 0.789389
R3423 VCC.n923 VCC.n922 0.789389
R3424 VCC.n924 VCC.n923 0.789389
R3425 VCC.n925 VCC.n924 0.789389
R3426 VCC.n926 VCC.n925 0.789389
R3427 VCC.n927 VCC.n926 0.789389
R3428 VCC.n928 VCC.n927 0.789389
R3429 VCC.n929 VCC.n928 0.789389
R3430 VCC.n930 VCC.n929 0.789389
R3431 VCC.n931 VCC.n930 0.789389
R3432 VCC.n1063 VCC.n1062 0.740931
R3433 VCC.n15 VCC.n14 0.6255
R3434 VCC.n1035 VCC.n1034 0.570812
R3435 VCC.n1037 VCC.n1036 0.570812
R3436 VCC.n1034 VCC.n1033 0.563
R3437 VCC.n1039 VCC.n1035 0.555188
R3438 VCC.n1038 VCC.n1037 0.555188
R3439 VCC.n1032 VCC.n1031 0.533
R3440 VCC.n1049 VCC.n6 0.436595
R3441 VCC.n1042 VCC.n1040 0.352137
R3442 VCC.n1062 VCC.n1060 0.313756
R3443 VCC.n1035 VCC.n428 0.2755
R3444 VCC.n1040 VCC.n1039 0.272875
R3445 VCC.n1039 VCC.n227 0.2505
R3446 VCC.n1034 VCC.n629 0.2505
R3447 VCC.n1033 VCC.n830 0.2505
R3448 VCC.n1063 VCC.n1058 0.152698
R3449 VCC.n1055 VCC.n1054 0.102063
R3450 VCC.n1043 VCC.n1042 0.0223101
R3451 VCC.n1040 VCC.n26 0.00150007
R3452 VCC.n1058 VCC.n1056 0.00120336
R3453 VCC.n1062 VCC.n1061 0.00120336
R3454 VCC.n9 VCC.n8 0.00101448
R3455 VCC.n1047 VCC.n1046 0.00100742
R3456 VCC.n1053 VCC.n1050 0.00100741
R3457 VCC.n26 VCC.n25 0.00100167
R3458 VCC.n17 VCC.n16 0.00100027
R3459 VCC.n19 VCC.n18 0.00100007
R3460 VCC.n1043 VCC.n10 0.00100006
R3461 VCC.n1049 VCC.n1043 0.00100001
R3462 VCC.n1050 VCC.n1049 0.001
R3463 VCC.n1033 VCC.n1032 0.001
R3464 VCC.n1049 VCC.n9 0.001
R3465 VCC.n1049 VCC.n1047 0.001
R3466 VCC.n1049 VCC.n1048 0.001
R3467 VCC.n1054 VCC.n5 0.000548326
R3468 VCC.n1042 VCC.n1041 0.000548326
R3469 VCC.n1054 VCC.n4 0.000548326
R3470 VCC.n1054 VCC.n1053 0.000548326
R3471 VCC.n1046 VCC.n1045 0.000507061
R3472 VCC.n4 VCC.n3 0.000507061
R3473 VCC.n3 VCC.n2 0.000507061
R3474 VCC.n1053 VCC.n1052 0.000507061
R3475 VCC.n2 VCC.n1 0.000507061
R3476 VCC.n15 VCC.n17 0.000500289
R3477 VCC.n22 VCC.n21 0.000500185
R3478 VCC.n12 VCC.n11 0.000500108
R3479 VCC.n13 VCC.n12 0.000500108
R3480 VCC.n20 VCC.n19 0.000500071
R3481 VCC.n1039 VCC.n1038 0.000500002
R3482 m9m10 m9m10.n498 25.8836
R3483 m9m10.n198 m9m10.n98 6.78175
R3484 m9m10.n513 m9m10.t511 6.70615
R3485 m9m10.n499 m9m10.t502 6.66895
R3486 m9m10.n99 m9m10.t423 6.50308
R3487 m9m10.n399 m9m10.t372 6.50308
R3488 m9m10.n299 m9m10.t386 6.50308
R3489 m9m10.n199 m9m10.t404 6.50308
R3490 m9m10.n0 m9m10.t29 6.50308
R3491 m9m10.n527 m9m10.n526 6.18831
R3492 m9m10.n109 m9m10.t368 5.71419
R3493 m9m10.n108 m9m10.t479 5.71419
R3494 m9m10.n107 m9m10.t111 5.71419
R3495 m9m10.n106 m9m10.t488 5.71419
R3496 m9m10.n105 m9m10.t325 5.71419
R3497 m9m10.n104 m9m10.t92 5.71419
R3498 m9m10.n103 m9m10.t301 5.71419
R3499 m9m10.n102 m9m10.t436 5.71419
R3500 m9m10.n101 m9m10.t207 5.71419
R3501 m9m10.n100 m9m10.t411 5.71419
R3502 m9m10.n99 m9m10.t193 5.71419
R3503 m9m10.n111 m9m10.t360 5.71419
R3504 m9m10.n112 m9m10.t120 5.71419
R3505 m9m10.n113 m9m10.t376 5.71419
R3506 m9m10.n114 m9m10.t50 5.71419
R3507 m9m10.n115 m9m10.t160 5.71419
R3508 m9m10.n116 m9m10.t44 5.71419
R3509 m9m10.n117 m9m10.t252 5.71419
R3510 m9m10.n118 m9m10.t62 5.71419
R3511 m9m10.n119 m9m10.t430 5.71419
R3512 m9m10.n120 m9m10.t171 5.71419
R3513 m9m10.n121 m9m10.t422 5.71419
R3514 m9m10.n122 m9m10.t452 5.71419
R3515 m9m10.n123 m9m10.t320 5.71419
R3516 m9m10.n124 m9m10.t106 5.71419
R3517 m9m10.n125 m9m10.t311 5.71419
R3518 m9m10.n126 m9m10.t121 5.71419
R3519 m9m10.n127 m9m10.t330 5.71419
R3520 m9m10.n128 m9m10.t221 5.71419
R3521 m9m10.n129 m9m10.t487 5.71419
R3522 m9m10.n130 m9m10.t61 5.71419
R3523 m9m10.n131 m9m10.t428 5.71419
R3524 m9m10.n132 m9m10.t54 5.71419
R3525 m9m10.n133 m9m10.t417 5.71419
R3526 m9m10.n134 m9m10.t288 5.71419
R3527 m9m10.n135 m9m10.t444 5.71419
R3528 m9m10.n136 m9m10.t309 5.71419
R3529 m9m10.n137 m9m10.t66 5.71419
R3530 m9m10.n138 m9m10.t298 5.71419
R3531 m9m10.n139 m9m10.t494 5.71419
R3532 m9m10.n140 m9m10.t115 5.71419
R3533 m9m10.n141 m9m10.t485 5.71419
R3534 m9m10.n142 m9m10.t215 5.71419
R3535 m9m10.n143 m9m10.t4 5.71419
R3536 m9m10.n144 m9m10.t365 5.71419
R3537 m9m10.n145 m9m10.t124 5.71419
R3538 m9m10.n146 m9m10.t359 5.71419
R3539 m9m10.n147 m9m10.t382 5.71419
R3540 m9m10.n148 m9m10.t265 5.71419
R3541 m9m10.n149 m9m10.t48 5.71419
R3542 m9m10.n150 m9m10.t256 5.71419
R3543 m9m10.n151 m9m10.t67 5.71419
R3544 m9m10.n152 m9m10.t275 5.71419
R3545 m9m10.n153 m9m10.t175 5.71419
R3546 m9m10.n154 m9m10.t427 5.71419
R3547 m9m10.n155 m9m10.t425 5.71419
R3548 m9m10.n156 m9m10.t324 5.71419
R3549 m9m10.n157 m9m10.t448 5.71419
R3550 m9m10.n158 m9m10.t316 5.71419
R3551 m9m10.n159 m9m10.t212 5.71419
R3552 m9m10.n160 m9m10.t334 5.71419
R3553 m9m10.n161 m9m10.t225 5.71419
R3554 m9m10.n162 m9m10.t460 5.71419
R3555 m9m10.n163 m9m10.t492 5.71419
R3556 m9m10.n164 m9m10.t375 5.71419
R3557 m9m10.n165 m9m10.t9 5.71419
R3558 m9m10.n166 m9m10.t370 5.71419
R3559 m9m10.n167 m9m10.t129 5.71419
R3560 m9m10.n168 m9m10.t387 5.71419
R3561 m9m10.n169 m9m10.t273 5.71419
R3562 m9m10.n170 m9m10.t20 5.71419
R3563 m9m10.n171 m9m10.t56 5.71419
R3564 m9m10.n172 m9m10.t261 5.71419
R3565 m9m10.n173 m9m10.t188 5.71419
R3566 m9m10.n174 m9m10.t445 5.71419
R3567 m9m10.n175 m9m10.t180 5.71419
R3568 m9m10.n176 m9m10.t434 5.71419
R3569 m9m10.n177 m9m10.t201 5.71419
R3570 m9m10.n178 m9m10.t86 5.71419
R3571 m9m10.n179 m9m10.t117 5.71419
R3572 m9m10.n180 m9m10.t322 5.71419
R3573 m9m10.n181 m9m10.t234 5.71419
R3574 m9m10.n182 m9m10.t338 5.71419
R3575 m9m10.n183 m9m10.t229 5.71419
R3576 m9m10.n184 m9m10.t125 5.71419
R3577 m9m10.n185 m9m10.t241 5.71419
R3578 m9m10.n186 m9m10.t141 5.71419
R3579 m9m10.n187 m9m10.t139 5.71419
R3580 m9m10.n188 m9m10.t374 5.71419
R3581 m9m10.n189 m9m10.t259 5.71419
R3582 m9m10.n190 m9m10.t395 5.71419
R3583 m9m10.n191 m9m10.t276 5.71419
R3584 m9m10.n192 m9m10.t26 5.71419
R3585 m9m10.n193 m9m10.t270 5.71419
R3586 m9m10.n194 m9m10.t196 5.71419
R3587 m9m10.n195 m9m10.t192 5.71419
R3588 m9m10.n196 m9m10.t450 5.71419
R3589 m9m10.n197 m9m10.t186 5.71419
R3590 m9m10.n497 m9m10.t294 5.71419
R3591 m9m10.n496 m9m10.t97 5.71419
R3592 m9m10.n495 m9m10.t305 5.71419
R3593 m9m10.n494 m9m10.t307 5.71419
R3594 m9m10.n493 m9m10.t406 5.71419
R3595 m9m10.n492 m9m10.t161 5.71419
R3596 m9m10.n491 m9m10.t416 5.71419
R3597 m9m10.n490 m9m10.t53 5.71419
R3598 m9m10.n489 m9m10.t390 5.71419
R3599 m9m10.n488 m9m10.t30 5.71419
R3600 m9m10.n487 m9m10.t248 5.71419
R3601 m9m10.n486 m9m10.t250 5.71419
R3602 m9m10.n485 m9m10.t369 5.71419
R3603 m9m10.n484 m9m10.t238 5.71419
R3604 m9m10.n483 m9m10.t350 5.71419
R3605 m9m10.n482 m9m10.t489 5.71419
R3606 m9m10.n481 m9m10.t357 5.71419
R3607 m9m10.n480 m9m10.t466 5.71419
R3608 m9m10.n479 m9m10.t232 5.71419
R3609 m9m10.n478 m9m10.t210 5.71419
R3610 m9m10.n477 m9m10.t312 5.71419
R3611 m9m10.n476 m9m10.t79 5.71419
R3612 m9m10.n475 m9m10.t291 5.71419
R3613 m9m10.n474 m9m10.t89 5.71419
R3614 m9m10.n473 m9m10.t296 5.71419
R3615 m9m10.n472 m9m10.t396 5.71419
R3616 m9m10.n471 m9m10.t185 5.71419
R3617 m9m10.n470 m9m10.t156 5.71419
R3618 m9m10.n469 m9m10.t408 5.71419
R3619 m9m10.n468 m9m10.t46 5.71419
R3620 m9m10.n467 m9m10.t242 5.71419
R3621 m9m10.n466 m9m10.t23 5.71419
R3622 m9m10.n465 m9m10.t146 5.71419
R3623 m9m10.n464 m9m10.t32 5.71419
R3624 m9m10.n463 m9m10.t132 5.71419
R3625 m9m10.n462 m9m10.t107 5.71419
R3626 m9m10.n461 m9m10.t344 5.71419
R3627 m9m10.n460 m9m10.t480 5.71419
R3628 m9m10.n459 m9m10.t331 5.71419
R3629 m9m10.n458 m9m10.t462 5.71419
R3630 m9m10.n457 m9m10.t95 5.71419
R3631 m9m10.n456 m9m10.t467 5.71419
R3632 m9m10.n455 m9m10.t73 5.71419
R3633 m9m10.n454 m9m10.t74 5.71419
R3634 m9m10.n453 m9m10.t286 5.71419
R3635 m9m10.n452 m9m10.t414 5.71419
R3636 m9m10.n451 m9m10.t198 5.71419
R3637 m9m10.n450 m9m10.t388 5.71419
R3638 m9m10.n449 m9m10.t176 5.71419
R3639 m9m10.n448 m9m10.t397 5.71419
R3640 m9m10.n447 m9m10.t37 5.71419
R3641 m9m10.n446 m9m10.t10 5.71419
R3642 m9m10.n445 m9m10.t237 5.71419
R3643 m9m10.n444 m9m10.t15 5.71419
R3644 m9m10.n443 m9m10.t143 5.71419
R3645 m9m10.n442 m9m10.t335 5.71419
R3646 m9m10.n441 m9m10.t126 5.71419
R3647 m9m10.n440 m9m10.t231 5.71419
R3648 m9m10.n439 m9m10.t133 5.71419
R3649 m9m10.n438 m9m10.t451 5.71419
R3650 m9m10.n437 m9m10.t194 5.71419
R3651 m9m10.n436 m9m10.t456 5.71419
R3652 m9m10.n435 m9m10.t87 5.71419
R3653 m9m10.n434 m9m10.t439 5.71419
R3654 m9m10.n433 m9m10.t68 5.71419
R3655 m9m10.n432 m9m10.t184 5.71419
R3656 m9m10.n431 m9m10.t75 5.71419
R3657 m9m10.n430 m9m10.t189 5.71419
R3658 m9m10.n429 m9m10.t446 5.71419
R3659 m9m10.n428 m9m10.t191 5.71419
R3660 m9m10.n427 m9m10.t287 5.71419
R3661 m9m10.n426 m9m10.t84 5.71419
R3662 m9m10.n425 m9m10.t274 5.71419
R3663 m9m10.n424 m9m10.t64 5.71419
R3664 m9m10.n423 m9m10.t278 5.71419
R3665 m9m10.n422 m9m10.t400 5.71419
R3666 m9m10.n421 m9m10.t371 5.71419
R3667 m9m10.n420 m9m10.t136 5.71419
R3668 m9m10.n419 m9m10.t380 5.71419
R3669 m9m10.n418 m9m10.t17 5.71419
R3670 m9m10.n417 m9m10.t226 5.71419
R3671 m9m10.n416 m9m10.t1 5.71419
R3672 m9m10.n415 m9m10.t127 5.71419
R3673 m9m10.n414 m9m10.t8 5.71419
R3674 m9m10.n413 m9m10.t340 5.71419
R3675 m9m10.n412 m9m10.t81 5.71419
R3676 m9m10.n411 m9m10.t327 5.71419
R3677 m9m10.n410 m9m10.t457 5.71419
R3678 m9m10.n409 m9m10.t333 5.71419
R3679 m9m10.n408 m9m10.t441 5.71419
R3680 m9m10.n407 m9m10.t69 5.71419
R3681 m9m10.n406 m9m10.t447 5.71419
R3682 m9m10.n405 m9m10.t281 5.71419
R3683 m9m10.n404 m9m10.t52 5.71419
R3684 m9m10.n403 m9m10.t267 5.71419
R3685 m9m10.n402 m9m10.t383 5.71419
R3686 m9m10.n401 m9m10.t173 5.71419
R3687 m9m10.n400 m9m10.t367 5.71419
R3688 m9m10.n399 m9m10.t158 5.71419
R3689 m9m10.n397 m9m10.t253 5.71419
R3690 m9m10.n396 m9m10.t47 5.71419
R3691 m9m10.n395 m9m10.t262 5.71419
R3692 m9m10.n394 m9m10.t264 5.71419
R3693 m9m10.n393 m9m10.t355 5.71419
R3694 m9m10.n392 m9m10.t122 5.71419
R3695 m9m10.n391 m9m10.t363 5.71419
R3696 m9m10.n390 m9m10.t2 5.71419
R3697 m9m10.n389 m9m10.t346 5.71419
R3698 m9m10.n388 m9m10.t482 5.71419
R3699 m9m10.n387 m9m10.t218 5.71419
R3700 m9m10.n386 m9m10.t220 5.71419
R3701 m9m10.n385 m9m10.t328 5.71419
R3702 m9m10.n384 m9m10.t205 5.71419
R3703 m9m10.n383 m9m10.t306 5.71419
R3704 m9m10.n382 m9m10.t442 5.71419
R3705 m9m10.n381 m9m10.t317 5.71419
R3706 m9m10.n380 m9m10.t415 5.71419
R3707 m9m10.n379 m9m10.t199 5.71419
R3708 m9m10.n378 m9m10.t169 5.71419
R3709 m9m10.n377 m9m10.t268 5.71419
R3710 m9m10.n376 m9m10.t31 5.71419
R3711 m9m10.n375 m9m10.t249 5.71419
R3712 m9m10.n374 m9m10.t41 5.71419
R3713 m9m10.n373 m9m10.t257 5.71419
R3714 m9m10.n372 m9m10.t349 5.71419
R3715 m9m10.n371 m9m10.t144 5.71419
R3716 m9m10.n370 m9m10.t118 5.71419
R3717 m9m10.n369 m9m10.t358 5.71419
R3718 m9m10.n368 m9m10.t497 5.71419
R3719 m9m10.n367 m9m10.t209 5.71419
R3720 m9m10.n366 m9m10.t475 5.71419
R3721 m9m10.n365 m9m10.t108 5.71419
R3722 m9m10.n364 m9m10.t484 5.71419
R3723 m9m10.n363 m9m10.t88 5.71419
R3724 m9m10.n362 m9m10.t58 5.71419
R3725 m9m10.n361 m9m10.t297 5.71419
R3726 m9m10.n360 m9m10.t431 5.71419
R3727 m9m10.n359 m9m10.t280 5.71419
R3728 m9m10.n358 m9m10.t407 5.71419
R3729 m9m10.n357 m9m10.t45 5.71419
R3730 m9m10.n356 m9m10.t418 5.71419
R3731 m9m10.n355 m9m10.t22 5.71419
R3732 m9m10.n354 m9m10.t24 5.71419
R3733 m9m10.n353 m9m10.t246 5.71419
R3734 m9m10.n352 m9m10.t361 5.71419
R3735 m9m10.n351 m9m10.t153 5.71419
R3736 m9m10.n350 m9m10.t343 5.71419
R3737 m9m10.n349 m9m10.t135 5.71419
R3738 m9m10.n348 m9m10.t351 5.71419
R3739 m9m10.n347 m9m10.t490 5.71419
R3740 m9m10.n346 m9m10.t463 5.71419
R3741 m9m10.n345 m9m10.t204 5.71419
R3742 m9m10.n344 m9m10.t469 5.71419
R3743 m9m10.n343 m9m10.t103 5.71419
R3744 m9m10.n342 m9m10.t285 5.71419
R3745 m9m10.n341 m9m10.t80 5.71419
R3746 m9m10.n340 m9m10.t197 5.71419
R3747 m9m10.n339 m9m10.t91 5.71419
R3748 m9m10.n338 m9m10.t389 5.71419
R3749 m9m10.n337 m9m10.t151 5.71419
R3750 m9m10.n336 m9m10.t398 5.71419
R3751 m9m10.n335 m9m10.t38 5.71419
R3752 m9m10.n334 m9m10.t377 5.71419
R3753 m9m10.n333 m9m10.t14 5.71419
R3754 m9m10.n332 m9m10.t142 5.71419
R3755 m9m10.n331 m9m10.t25 5.71419
R3756 m9m10.n330 m9m10.t148 5.71419
R3757 m9m10.n329 m9m10.t459 5.71419
R3758 m9m10.n328 m9m10.t203 5.71419
R3759 m9m10.n327 m9m10.t300 5.71419
R3760 m9m10.n326 m9m10.t101 5.71419
R3761 m9m10.n325 m9m10.t282 5.71419
R3762 m9m10.n324 m9m10.t77 5.71419
R3763 m9m10.n323 m9m10.t290 5.71419
R3764 m9m10.n322 m9m10.t421 5.71419
R3765 m9m10.n321 m9m10.t385 5.71419
R3766 m9m10.n320 m9m10.t149 5.71419
R3767 m9m10.n319 m9m10.t394 5.71419
R3768 m9m10.n318 m9m10.t34 5.71419
R3769 m9m10.n317 m9m10.t235 5.71419
R3770 m9m10.n316 m9m10.t12 5.71419
R3771 m9m10.n315 m9m10.t137 5.71419
R3772 m9m10.n314 m9m10.t21 5.71419
R3773 m9m10.n313 m9m10.t353 5.71419
R3774 m9m10.n312 m9m10.t98 5.71419
R3775 m9m10.n311 m9m10.t337 5.71419
R3776 m9m10.n310 m9m10.t470 5.71419
R3777 m9m10.n309 m9m10.t342 5.71419
R3778 m9m10.n308 m9m10.t453 5.71419
R3779 m9m10.n307 m9m10.t82 5.71419
R3780 m9m10.n306 m9m10.t461 5.71419
R3781 m9m10.n305 m9m10.t292 5.71419
R3782 m9m10.n304 m9m10.t65 5.71419
R3783 m9m10.n303 m9m10.t277 5.71419
R3784 m9m10.n302 m9m10.t399 5.71419
R3785 m9m10.n301 m9m10.t187 5.71419
R3786 m9m10.n300 m9m10.t378 5.71419
R3787 m9m10.n299 m9m10.t170 5.71419
R3788 m9m10.n297 m9m10.t222 5.71419
R3789 m9m10.n296 m9m10.t498 5.71419
R3790 m9m10.n295 m9m10.t228 5.71419
R3791 m9m10.n294 m9m10.t230 5.71419
R3792 m9m10.n293 m9m10.t314 5.71419
R3793 m9m10.n292 m9m10.t76 5.71419
R3794 m9m10.n291 m9m10.t323 5.71419
R3795 m9m10.n290 m9m10.t455 5.71419
R3796 m9m10.n289 m9m10.t299 5.71419
R3797 m9m10.n288 m9m10.t433 5.71419
R3798 m9m10.n287 m9m10.t179 5.71419
R3799 m9m10.n286 m9m10.t182 5.71419
R3800 m9m10.n285 m9m10.t279 5.71419
R3801 m9m10.n284 m9m10.t166 5.71419
R3802 m9m10.n283 m9m10.t263 5.71419
R3803 m9m10.n282 m9m10.t381 5.71419
R3804 m9m10.n281 m9m10.t271 5.71419
R3805 m9m10.n280 m9m10.t362 5.71419
R3806 m9m10.n279 m9m10.t154 5.71419
R3807 m9m10.n278 m9m10.t130 5.71419
R3808 m9m10.n277 m9m10.t233 5.71419
R3809 m9m10.n276 m9m10.t483 5.71419
R3810 m9m10.n275 m9m10.t219 5.71419
R3811 m9m10.n274 m9m10.t493 5.71419
R3812 m9m10.n273 m9m10.t224 5.71419
R3813 m9m10.n272 m9m10.t304 5.71419
R3814 m9m10.n271 m9m10.t104 5.71419
R3815 m9m10.n270 m9m10.t71 5.71419
R3816 m9m10.n269 m9m10.t318 5.71419
R3817 m9m10.n268 m9m10.t449 5.71419
R3818 m9m10.n267 m9m10.t168 5.71419
R3819 m9m10.n266 m9m10.t426 5.71419
R3820 m9m10.n265 m9m10.t60 5.71419
R3821 m9m10.n264 m9m10.t435 5.71419
R3822 m9m10.n263 m9m10.t40 5.71419
R3823 m9m10.n262 m9m10.t6 5.71419
R3824 m9m10.n261 m9m10.t258 5.71419
R3825 m9m10.n260 m9m10.t373 5.71419
R3826 m9m10.n259 m9m10.t243 5.71419
R3827 m9m10.n258 m9m10.t356 5.71419
R3828 m9m10.n257 m9m10.t496 5.71419
R3829 m9m10.n256 m9m10.t364 5.71419
R3830 m9m10.n255 m9m10.t474 5.71419
R3831 m9m10.n254 m9m10.t476 5.71419
R3832 m9m10.n253 m9m10.t216 5.71419
R3833 m9m10.n252 m9m10.t321 5.71419
R3834 m9m10.n251 m9m10.t116 5.71419
R3835 m9m10.n250 m9m10.t295 5.71419
R3836 m9m10.n249 m9m10.t99 5.71419
R3837 m9m10.n248 m9m10.t308 5.71419
R3838 m9m10.n247 m9m10.t443 5.71419
R3839 m9m10.n246 m9m10.t409 5.71419
R3840 m9m10.n245 m9m10.t164 5.71419
R3841 m9m10.n244 m9m10.t419 5.71419
R3842 m9m10.n243 m9m10.t55 5.71419
R3843 m9m10.n242 m9m10.t245 5.71419
R3844 m9m10.n241 m9m10.t33 5.71419
R3845 m9m10.n240 m9m10.t152 5.71419
R3846 m9m10.n239 m9m10.t42 5.71419
R3847 m9m10.n238 m9m10.t345 5.71419
R3848 m9m10.n237 m9m10.t114 5.71419
R3849 m9m10.n236 m9m10.t352 5.71419
R3850 m9m10.n235 m9m10.t491 5.71419
R3851 m9m10.n234 m9m10.t336 5.71419
R3852 m9m10.n233 m9m10.t468 5.71419
R3853 m9m10.n232 m9m10.t102 5.71419
R3854 m9m10.n231 m9m10.t477 5.71419
R3855 m9m10.n230 m9m10.t109 5.71419
R3856 m9m10.n229 m9m10.t471 5.71419
R3857 m9m10.n228 m9m10.t213 5.71419
R3858 m9m10.n227 m9m10.t319 5.71419
R3859 m9m10.n226 m9m10.t112 5.71419
R3860 m9m10.n225 m9m10.t293 5.71419
R3861 m9m10.n224 m9m10.t93 5.71419
R3862 m9m10.n223 m9m10.t302 5.71419
R3863 m9m10.n222 m9m10.t437 5.71419
R3864 m9m10.n221 m9m10.t402 5.71419
R3865 m9m10.n220 m9m10.t159 5.71419
R3866 m9m10.n219 m9m10.t413 5.71419
R3867 m9m10.n218 m9m10.t49 5.71419
R3868 m9m10.n217 m9m10.t244 5.71419
R3869 m9m10.n216 m9m10.t27 5.71419
R3870 m9m10.n215 m9m10.t150 5.71419
R3871 m9m10.n214 m9m10.t35 5.71419
R3872 m9m10.n213 m9m10.t366 5.71419
R3873 m9m10.n212 m9m10.t110 5.71419
R3874 m9m10.n211 m9m10.t348 5.71419
R3875 m9m10.n210 m9m10.t486 5.71419
R3876 m9m10.n209 m9m10.t354 5.71419
R3877 m9m10.n208 m9m10.t464 5.71419
R3878 m9m10.n207 m9m10.t100 5.71419
R3879 m9m10.n206 m9m10.t472 5.71419
R3880 m9m10.n205 m9m10.t310 5.71419
R3881 m9m10.n204 m9m10.t78 5.71419
R3882 m9m10.n203 m9m10.t289 5.71419
R3883 m9m10.n202 m9m10.t420 5.71419
R3884 m9m10.n201 m9m10.t202 5.71419
R3885 m9m10.n200 m9m10.t392 5.71419
R3886 m9m10.n199 m9m10.t181 5.71419
R3887 m9m10.n98 m9m10.t391 5.71419
R3888 m9m10.n97 m9m10.t178 5.71419
R3889 m9m10.n96 m9m10.t401 5.71419
R3890 m9m10.n95 m9m10.t403 5.71419
R3891 m9m10.n94 m9m10.t11 5.71419
R3892 m9m10.n93 m9m10.t239 5.71419
R3893 m9m10.n92 m9m10.t18 5.71419
R3894 m9m10.n91 m9m10.t145 5.71419
R3895 m9m10.n90 m9m10.t3 5.71419
R3896 m9m10.n89 m9m10.t128 5.71419
R3897 m9m10.n88 m9m10.t339 5.71419
R3898 m9m10.n87 m9m10.t341 5.71419
R3899 m9m10.n86 m9m10.t478 5.71419
R3900 m9m10.n85 m9m10.t329 5.71419
R3901 m9m10.n84 m9m10.t458 5.71419
R3902 m9m10.n83 m9m10.t90 5.71419
R3903 m9m10.n82 m9m10.t465 5.71419
R3904 m9m10.n81 m9m10.t70 5.71419
R3905 m9m10.n80 m9m10.t315 5.71419
R3906 m9m10.n79 m9m10.t283 5.71419
R3907 m9m10.n78 m9m10.t410 5.71419
R3908 m9m10.n77 m9m10.t167 5.71419
R3909 m9m10.n76 m9m10.t384 5.71419
R3910 m9m10.n75 m9m10.t174 5.71419
R3911 m9m10.n74 m9m10.t393 5.71419
R3912 m9m10.n73 m9m10.t5 5.71419
R3913 m9m10.n72 m9m10.t255 5.71419
R3914 m9m10.n71 m9m10.t236 5.71419
R3915 m9m10.n70 m9m10.t13 5.71419
R3916 m9m10.n69 m9m10.t138 5.71419
R3917 m9m10.n68 m9m10.t332 5.71419
R3918 m9m10.n67 m9m10.t123 5.71419
R3919 m9m10.n66 m9m10.t227 5.71419
R3920 m9m10.n65 m9m10.t131 5.71419
R3921 m9m10.n64 m9m10.t214 5.71419
R3922 m9m10.n63 m9m10.t190 5.71419
R3923 m9m10.n62 m9m10.t454 5.71419
R3924 m9m10.n61 m9m10.t83 5.71419
R3925 m9m10.n60 m9m10.t432 5.71419
R3926 m9m10.n59 m9m10.t63 5.71419
R3927 m9m10.n58 m9m10.t177 5.71419
R3928 m9m10.n57 m9m10.t72 5.71419
R3929 m9m10.n56 m9m10.t162 5.71419
R3930 m9m10.n55 m9m10.t163 5.71419
R3931 m9m10.n54 m9m10.t379 5.71419
R3932 m9m10.n53 m9m10.t16 5.71419
R3933 m9m10.n52 m9m10.t269 5.71419
R3934 m9m10.n51 m9m10.t0 5.71419
R3935 m9m10.n50 m9m10.t251 5.71419
R3936 m9m10.n49 m9m10.t7 5.71419
R3937 m9m10.n48 m9m10.t134 5.71419
R3938 m9m10.n47 m9m10.t113 5.71419
R3939 m9m10.n46 m9m10.t326 5.71419
R3940 m9m10.n45 m9m10.t119 5.71419
R3941 m9m10.n44 m9m10.t223 5.71419
R3942 m9m10.n43 m9m10.t440 5.71419
R3943 m9m10.n42 m9m10.t211 5.71419
R3944 m9m10.n41 m9m10.t313 5.71419
R3945 m9m10.n40 m9m10.t217 5.71419
R3946 m9m10.n39 m9m10.t51 5.71419
R3947 m9m10.n38 m9m10.t266 5.71419
R3948 m9m10.n37 m9m10.t59 5.71419
R3949 m9m10.n36 m9m10.t172 5.71419
R3950 m9m10.n35 m9m10.t39 5.71419
R3951 m9m10.n34 m9m10.t157 5.71419
R3952 m9m10.n33 m9m10.t254 5.71419
R3953 m9m10.n32 m9m10.t165 5.71419
R3954 m9m10.n31 m9m10.t260 5.71419
R3955 m9m10.n30 m9m10.t94 5.71419
R3956 m9m10.n29 m9m10.t303 5.71419
R3957 m9m10.n28 m9m10.t438 5.71419
R3958 m9m10.n27 m9m10.t208 5.71419
R3959 m9m10.n26 m9m10.t412 5.71419
R3960 m9m10.n25 m9m10.t195 5.71419
R3961 m9m10.n24 m9m10.t424 5.71419
R3962 m9m10.n23 m9m10.t57 5.71419
R3963 m9m10.n22 m9m10.t28 5.71419
R3964 m9m10.n21 m9m10.t247 5.71419
R3965 m9m10.n20 m9m10.t36 5.71419
R3966 m9m10.n19 m9m10.t155 5.71419
R3967 m9m10.n18 m9m10.t347 5.71419
R3968 m9m10.n17 m9m10.t140 5.71419
R3969 m9m10.n16 m9m10.t240 5.71419
R3970 m9m10.n15 m9m10.t147 5.71419
R3971 m9m10.n14 m9m10.t495 5.71419
R3972 m9m10.n13 m9m10.t206 5.71419
R3973 m9m10.n12 m9m10.t473 5.71419
R3974 m9m10.n11 m9m10.t105 5.71419
R3975 m9m10.n10 m9m10.t481 5.71419
R3976 m9m10.n9 m9m10.t85 5.71419
R3977 m9m10.n8 m9m10.t200 5.71419
R3978 m9m10.n7 m9m10.t96 5.71419
R3979 m9m10.n6 m9m10.t429 5.71419
R3980 m9m10.n5 m9m10.t183 5.71419
R3981 m9m10.n4 m9m10.t405 5.71419
R3982 m9m10.n3 m9m10.t43 5.71419
R3983 m9m10.n2 m9m10.t284 5.71419
R3984 m9m10.n1 m9m10.t19 5.71419
R3985 m9m10.n0 m9m10.t272 5.71419
R3986 m9m10.n512 m9m10.t500 5.71419
R3987 m9m10.n511 m9m10.t527 5.71419
R3988 m9m10.n510 m9m10.t526 5.71419
R3989 m9m10.n509 m9m10.t522 5.71419
R3990 m9m10.n508 m9m10.t513 5.71419
R3991 m9m10.n507 m9m10.t504 5.71419
R3992 m9m10.n506 m9m10.t510 5.71419
R3993 m9m10.n505 m9m10.t525 5.71419
R3994 m9m10.n504 m9m10.t512 5.71419
R3995 m9m10.n503 m9m10.t523 5.71419
R3996 m9m10.n502 m9m10.t519 5.71419
R3997 m9m10.n501 m9m10.t514 5.71419
R3998 m9m10.n500 m9m10.t503 5.71419
R3999 m9m10.n499 m9m10.t517 5.71419
R4000 m9m10.n526 m9m10.t509 5.71419
R4001 m9m10.n525 m9m10.t516 5.71419
R4002 m9m10.n524 m9m10.t507 5.71419
R4003 m9m10.n523 m9m10.t506 5.71419
R4004 m9m10.n522 m9m10.t521 5.71419
R4005 m9m10.n521 m9m10.t524 5.71419
R4006 m9m10.n520 m9m10.t518 5.71419
R4007 m9m10.n519 m9m10.t505 5.71419
R4008 m9m10.n518 m9m10.t520 5.71419
R4009 m9m10.n517 m9m10.t508 5.71419
R4010 m9m10.n516 m9m10.t501 5.71419
R4011 m9m10.n515 m9m10.t528 5.71419
R4012 m9m10.n514 m9m10.t515 5.71419
R4013 m9m10.n513 m9m10.t529 5.71419
R4014 m9m10.n110 m9m10.t499 5.71419
R4015 m9m10.n527 m9m10.n512 5.42983
R4016 m9m10.n298 m9m10.n198 4.5005
R4017 m9m10.n398 m9m10.n298 4.5005
R4018 m9m10.n498 m9m10.n398 4.5005
R4019 m9m10.n498 m9m10.n497 2.34425
R4020 m9m10.n398 m9m10.n397 2.34425
R4021 m9m10.n298 m9m10.n297 2.34425
R4022 m9m10.n198 m9m10.n197 2.34425
R4023 m9m10.n514 m9m10.n513 0.992464
R4024 m9m10.n515 m9m10.n514 0.992464
R4025 m9m10.n516 m9m10.n515 0.992464
R4026 m9m10.n517 m9m10.n516 0.992464
R4027 m9m10.n518 m9m10.n517 0.992464
R4028 m9m10.n519 m9m10.n518 0.992464
R4029 m9m10.n520 m9m10.n519 0.992464
R4030 m9m10.n521 m9m10.n520 0.992464
R4031 m9m10.n522 m9m10.n521 0.992464
R4032 m9m10.n523 m9m10.n522 0.992464
R4033 m9m10.n524 m9m10.n523 0.992464
R4034 m9m10.n525 m9m10.n524 0.992464
R4035 m9m10.n526 m9m10.n525 0.992464
R4036 m9m10.n500 m9m10.n499 0.955262
R4037 m9m10.n501 m9m10.n500 0.955262
R4038 m9m10.n502 m9m10.n501 0.955262
R4039 m9m10.n503 m9m10.n502 0.955262
R4040 m9m10.n504 m9m10.n503 0.955262
R4041 m9m10.n505 m9m10.n504 0.955262
R4042 m9m10.n506 m9m10.n505 0.955262
R4043 m9m10.n507 m9m10.n506 0.955262
R4044 m9m10.n508 m9m10.n507 0.955262
R4045 m9m10.n509 m9m10.n508 0.955262
R4046 m9m10.n510 m9m10.n509 0.955262
R4047 m9m10.n511 m9m10.n510 0.955262
R4048 m9m10.n512 m9m10.n511 0.955262
R4049 m9m10 m9m10.n527 0.8205
R4050 m9m10.n100 m9m10.n99 0.789389
R4051 m9m10.n101 m9m10.n100 0.789389
R4052 m9m10.n102 m9m10.n101 0.789389
R4053 m9m10.n103 m9m10.n102 0.789389
R4054 m9m10.n104 m9m10.n103 0.789389
R4055 m9m10.n105 m9m10.n104 0.789389
R4056 m9m10.n106 m9m10.n105 0.789389
R4057 m9m10.n107 m9m10.n106 0.789389
R4058 m9m10.n108 m9m10.n107 0.789389
R4059 m9m10.n109 m9m10.n108 0.789389
R4060 m9m10.n110 m9m10.n109 0.789389
R4061 m9m10.n400 m9m10.n399 0.789389
R4062 m9m10.n401 m9m10.n400 0.789389
R4063 m9m10.n402 m9m10.n401 0.789389
R4064 m9m10.n403 m9m10.n402 0.789389
R4065 m9m10.n404 m9m10.n403 0.789389
R4066 m9m10.n405 m9m10.n404 0.789389
R4067 m9m10.n406 m9m10.n405 0.789389
R4068 m9m10.n407 m9m10.n406 0.789389
R4069 m9m10.n408 m9m10.n407 0.789389
R4070 m9m10.n409 m9m10.n408 0.789389
R4071 m9m10.n410 m9m10.n409 0.789389
R4072 m9m10.n411 m9m10.n410 0.789389
R4073 m9m10.n412 m9m10.n411 0.789389
R4074 m9m10.n413 m9m10.n412 0.789389
R4075 m9m10.n414 m9m10.n413 0.789389
R4076 m9m10.n415 m9m10.n414 0.789389
R4077 m9m10.n416 m9m10.n415 0.789389
R4078 m9m10.n417 m9m10.n416 0.789389
R4079 m9m10.n418 m9m10.n417 0.789389
R4080 m9m10.n419 m9m10.n418 0.789389
R4081 m9m10.n420 m9m10.n419 0.789389
R4082 m9m10.n421 m9m10.n420 0.789389
R4083 m9m10.n422 m9m10.n421 0.789389
R4084 m9m10.n423 m9m10.n422 0.789389
R4085 m9m10.n424 m9m10.n423 0.789389
R4086 m9m10.n425 m9m10.n424 0.789389
R4087 m9m10.n426 m9m10.n425 0.789389
R4088 m9m10.n427 m9m10.n426 0.789389
R4089 m9m10.n428 m9m10.n427 0.789389
R4090 m9m10.n429 m9m10.n428 0.789389
R4091 m9m10.n430 m9m10.n429 0.789389
R4092 m9m10.n431 m9m10.n430 0.789389
R4093 m9m10.n432 m9m10.n431 0.789389
R4094 m9m10.n433 m9m10.n432 0.789389
R4095 m9m10.n434 m9m10.n433 0.789389
R4096 m9m10.n435 m9m10.n434 0.789389
R4097 m9m10.n436 m9m10.n435 0.789389
R4098 m9m10.n437 m9m10.n436 0.789389
R4099 m9m10.n438 m9m10.n437 0.789389
R4100 m9m10.n439 m9m10.n438 0.789389
R4101 m9m10.n440 m9m10.n439 0.789389
R4102 m9m10.n441 m9m10.n440 0.789389
R4103 m9m10.n442 m9m10.n441 0.789389
R4104 m9m10.n443 m9m10.n442 0.789389
R4105 m9m10.n444 m9m10.n443 0.789389
R4106 m9m10.n445 m9m10.n444 0.789389
R4107 m9m10.n446 m9m10.n445 0.789389
R4108 m9m10.n447 m9m10.n446 0.789389
R4109 m9m10.n448 m9m10.n447 0.789389
R4110 m9m10.n449 m9m10.n448 0.789389
R4111 m9m10.n450 m9m10.n449 0.789389
R4112 m9m10.n451 m9m10.n450 0.789389
R4113 m9m10.n452 m9m10.n451 0.789389
R4114 m9m10.n453 m9m10.n452 0.789389
R4115 m9m10.n454 m9m10.n453 0.789389
R4116 m9m10.n455 m9m10.n454 0.789389
R4117 m9m10.n456 m9m10.n455 0.789389
R4118 m9m10.n457 m9m10.n456 0.789389
R4119 m9m10.n458 m9m10.n457 0.789389
R4120 m9m10.n459 m9m10.n458 0.789389
R4121 m9m10.n460 m9m10.n459 0.789389
R4122 m9m10.n461 m9m10.n460 0.789389
R4123 m9m10.n462 m9m10.n461 0.789389
R4124 m9m10.n463 m9m10.n462 0.789389
R4125 m9m10.n464 m9m10.n463 0.789389
R4126 m9m10.n465 m9m10.n464 0.789389
R4127 m9m10.n466 m9m10.n465 0.789389
R4128 m9m10.n467 m9m10.n466 0.789389
R4129 m9m10.n468 m9m10.n467 0.789389
R4130 m9m10.n469 m9m10.n468 0.789389
R4131 m9m10.n470 m9m10.n469 0.789389
R4132 m9m10.n471 m9m10.n470 0.789389
R4133 m9m10.n472 m9m10.n471 0.789389
R4134 m9m10.n473 m9m10.n472 0.789389
R4135 m9m10.n474 m9m10.n473 0.789389
R4136 m9m10.n475 m9m10.n474 0.789389
R4137 m9m10.n476 m9m10.n475 0.789389
R4138 m9m10.n477 m9m10.n476 0.789389
R4139 m9m10.n478 m9m10.n477 0.789389
R4140 m9m10.n479 m9m10.n478 0.789389
R4141 m9m10.n480 m9m10.n479 0.789389
R4142 m9m10.n481 m9m10.n480 0.789389
R4143 m9m10.n482 m9m10.n481 0.789389
R4144 m9m10.n483 m9m10.n482 0.789389
R4145 m9m10.n484 m9m10.n483 0.789389
R4146 m9m10.n485 m9m10.n484 0.789389
R4147 m9m10.n486 m9m10.n485 0.789389
R4148 m9m10.n487 m9m10.n486 0.789389
R4149 m9m10.n488 m9m10.n487 0.789389
R4150 m9m10.n489 m9m10.n488 0.789389
R4151 m9m10.n490 m9m10.n489 0.789389
R4152 m9m10.n491 m9m10.n490 0.789389
R4153 m9m10.n492 m9m10.n491 0.789389
R4154 m9m10.n493 m9m10.n492 0.789389
R4155 m9m10.n494 m9m10.n493 0.789389
R4156 m9m10.n495 m9m10.n494 0.789389
R4157 m9m10.n496 m9m10.n495 0.789389
R4158 m9m10.n497 m9m10.n496 0.789389
R4159 m9m10.n300 m9m10.n299 0.789389
R4160 m9m10.n301 m9m10.n300 0.789389
R4161 m9m10.n302 m9m10.n301 0.789389
R4162 m9m10.n303 m9m10.n302 0.789389
R4163 m9m10.n304 m9m10.n303 0.789389
R4164 m9m10.n305 m9m10.n304 0.789389
R4165 m9m10.n306 m9m10.n305 0.789389
R4166 m9m10.n307 m9m10.n306 0.789389
R4167 m9m10.n308 m9m10.n307 0.789389
R4168 m9m10.n309 m9m10.n308 0.789389
R4169 m9m10.n310 m9m10.n309 0.789389
R4170 m9m10.n311 m9m10.n310 0.789389
R4171 m9m10.n312 m9m10.n311 0.789389
R4172 m9m10.n313 m9m10.n312 0.789389
R4173 m9m10.n314 m9m10.n313 0.789389
R4174 m9m10.n315 m9m10.n314 0.789389
R4175 m9m10.n316 m9m10.n315 0.789389
R4176 m9m10.n317 m9m10.n316 0.789389
R4177 m9m10.n318 m9m10.n317 0.789389
R4178 m9m10.n319 m9m10.n318 0.789389
R4179 m9m10.n320 m9m10.n319 0.789389
R4180 m9m10.n321 m9m10.n320 0.789389
R4181 m9m10.n322 m9m10.n321 0.789389
R4182 m9m10.n323 m9m10.n322 0.789389
R4183 m9m10.n324 m9m10.n323 0.789389
R4184 m9m10.n325 m9m10.n324 0.789389
R4185 m9m10.n326 m9m10.n325 0.789389
R4186 m9m10.n327 m9m10.n326 0.789389
R4187 m9m10.n328 m9m10.n327 0.789389
R4188 m9m10.n329 m9m10.n328 0.789389
R4189 m9m10.n330 m9m10.n329 0.789389
R4190 m9m10.n331 m9m10.n330 0.789389
R4191 m9m10.n332 m9m10.n331 0.789389
R4192 m9m10.n333 m9m10.n332 0.789389
R4193 m9m10.n334 m9m10.n333 0.789389
R4194 m9m10.n335 m9m10.n334 0.789389
R4195 m9m10.n336 m9m10.n335 0.789389
R4196 m9m10.n337 m9m10.n336 0.789389
R4197 m9m10.n338 m9m10.n337 0.789389
R4198 m9m10.n339 m9m10.n338 0.789389
R4199 m9m10.n340 m9m10.n339 0.789389
R4200 m9m10.n341 m9m10.n340 0.789389
R4201 m9m10.n342 m9m10.n341 0.789389
R4202 m9m10.n343 m9m10.n342 0.789389
R4203 m9m10.n344 m9m10.n343 0.789389
R4204 m9m10.n345 m9m10.n344 0.789389
R4205 m9m10.n346 m9m10.n345 0.789389
R4206 m9m10.n347 m9m10.n346 0.789389
R4207 m9m10.n348 m9m10.n347 0.789389
R4208 m9m10.n349 m9m10.n348 0.789389
R4209 m9m10.n350 m9m10.n349 0.789389
R4210 m9m10.n351 m9m10.n350 0.789389
R4211 m9m10.n352 m9m10.n351 0.789389
R4212 m9m10.n353 m9m10.n352 0.789389
R4213 m9m10.n354 m9m10.n353 0.789389
R4214 m9m10.n355 m9m10.n354 0.789389
R4215 m9m10.n356 m9m10.n355 0.789389
R4216 m9m10.n357 m9m10.n356 0.789389
R4217 m9m10.n358 m9m10.n357 0.789389
R4218 m9m10.n359 m9m10.n358 0.789389
R4219 m9m10.n360 m9m10.n359 0.789389
R4220 m9m10.n361 m9m10.n360 0.789389
R4221 m9m10.n362 m9m10.n361 0.789389
R4222 m9m10.n363 m9m10.n362 0.789389
R4223 m9m10.n364 m9m10.n363 0.789389
R4224 m9m10.n365 m9m10.n364 0.789389
R4225 m9m10.n366 m9m10.n365 0.789389
R4226 m9m10.n367 m9m10.n366 0.789389
R4227 m9m10.n368 m9m10.n367 0.789389
R4228 m9m10.n369 m9m10.n368 0.789389
R4229 m9m10.n370 m9m10.n369 0.789389
R4230 m9m10.n371 m9m10.n370 0.789389
R4231 m9m10.n372 m9m10.n371 0.789389
R4232 m9m10.n373 m9m10.n372 0.789389
R4233 m9m10.n374 m9m10.n373 0.789389
R4234 m9m10.n375 m9m10.n374 0.789389
R4235 m9m10.n376 m9m10.n375 0.789389
R4236 m9m10.n377 m9m10.n376 0.789389
R4237 m9m10.n378 m9m10.n377 0.789389
R4238 m9m10.n379 m9m10.n378 0.789389
R4239 m9m10.n380 m9m10.n379 0.789389
R4240 m9m10.n381 m9m10.n380 0.789389
R4241 m9m10.n382 m9m10.n381 0.789389
R4242 m9m10.n383 m9m10.n382 0.789389
R4243 m9m10.n384 m9m10.n383 0.789389
R4244 m9m10.n385 m9m10.n384 0.789389
R4245 m9m10.n386 m9m10.n385 0.789389
R4246 m9m10.n387 m9m10.n386 0.789389
R4247 m9m10.n388 m9m10.n387 0.789389
R4248 m9m10.n389 m9m10.n388 0.789389
R4249 m9m10.n390 m9m10.n389 0.789389
R4250 m9m10.n391 m9m10.n390 0.789389
R4251 m9m10.n392 m9m10.n391 0.789389
R4252 m9m10.n393 m9m10.n392 0.789389
R4253 m9m10.n394 m9m10.n393 0.789389
R4254 m9m10.n395 m9m10.n394 0.789389
R4255 m9m10.n396 m9m10.n395 0.789389
R4256 m9m10.n397 m9m10.n396 0.789389
R4257 m9m10.n200 m9m10.n199 0.789389
R4258 m9m10.n201 m9m10.n200 0.789389
R4259 m9m10.n202 m9m10.n201 0.789389
R4260 m9m10.n203 m9m10.n202 0.789389
R4261 m9m10.n204 m9m10.n203 0.789389
R4262 m9m10.n205 m9m10.n204 0.789389
R4263 m9m10.n206 m9m10.n205 0.789389
R4264 m9m10.n207 m9m10.n206 0.789389
R4265 m9m10.n208 m9m10.n207 0.789389
R4266 m9m10.n209 m9m10.n208 0.789389
R4267 m9m10.n210 m9m10.n209 0.789389
R4268 m9m10.n211 m9m10.n210 0.789389
R4269 m9m10.n212 m9m10.n211 0.789389
R4270 m9m10.n213 m9m10.n212 0.789389
R4271 m9m10.n214 m9m10.n213 0.789389
R4272 m9m10.n215 m9m10.n214 0.789389
R4273 m9m10.n216 m9m10.n215 0.789389
R4274 m9m10.n217 m9m10.n216 0.789389
R4275 m9m10.n218 m9m10.n217 0.789389
R4276 m9m10.n219 m9m10.n218 0.789389
R4277 m9m10.n220 m9m10.n219 0.789389
R4278 m9m10.n221 m9m10.n220 0.789389
R4279 m9m10.n222 m9m10.n221 0.789389
R4280 m9m10.n223 m9m10.n222 0.789389
R4281 m9m10.n224 m9m10.n223 0.789389
R4282 m9m10.n225 m9m10.n224 0.789389
R4283 m9m10.n226 m9m10.n225 0.789389
R4284 m9m10.n227 m9m10.n226 0.789389
R4285 m9m10.n228 m9m10.n227 0.789389
R4286 m9m10.n229 m9m10.n228 0.789389
R4287 m9m10.n230 m9m10.n229 0.789389
R4288 m9m10.n231 m9m10.n230 0.789389
R4289 m9m10.n232 m9m10.n231 0.789389
R4290 m9m10.n233 m9m10.n232 0.789389
R4291 m9m10.n234 m9m10.n233 0.789389
R4292 m9m10.n235 m9m10.n234 0.789389
R4293 m9m10.n236 m9m10.n235 0.789389
R4294 m9m10.n237 m9m10.n236 0.789389
R4295 m9m10.n238 m9m10.n237 0.789389
R4296 m9m10.n239 m9m10.n238 0.789389
R4297 m9m10.n240 m9m10.n239 0.789389
R4298 m9m10.n241 m9m10.n240 0.789389
R4299 m9m10.n242 m9m10.n241 0.789389
R4300 m9m10.n243 m9m10.n242 0.789389
R4301 m9m10.n244 m9m10.n243 0.789389
R4302 m9m10.n245 m9m10.n244 0.789389
R4303 m9m10.n246 m9m10.n245 0.789389
R4304 m9m10.n247 m9m10.n246 0.789389
R4305 m9m10.n248 m9m10.n247 0.789389
R4306 m9m10.n249 m9m10.n248 0.789389
R4307 m9m10.n250 m9m10.n249 0.789389
R4308 m9m10.n251 m9m10.n250 0.789389
R4309 m9m10.n252 m9m10.n251 0.789389
R4310 m9m10.n253 m9m10.n252 0.789389
R4311 m9m10.n254 m9m10.n253 0.789389
R4312 m9m10.n255 m9m10.n254 0.789389
R4313 m9m10.n256 m9m10.n255 0.789389
R4314 m9m10.n257 m9m10.n256 0.789389
R4315 m9m10.n258 m9m10.n257 0.789389
R4316 m9m10.n259 m9m10.n258 0.789389
R4317 m9m10.n260 m9m10.n259 0.789389
R4318 m9m10.n261 m9m10.n260 0.789389
R4319 m9m10.n262 m9m10.n261 0.789389
R4320 m9m10.n263 m9m10.n262 0.789389
R4321 m9m10.n264 m9m10.n263 0.789389
R4322 m9m10.n265 m9m10.n264 0.789389
R4323 m9m10.n266 m9m10.n265 0.789389
R4324 m9m10.n267 m9m10.n266 0.789389
R4325 m9m10.n268 m9m10.n267 0.789389
R4326 m9m10.n269 m9m10.n268 0.789389
R4327 m9m10.n270 m9m10.n269 0.789389
R4328 m9m10.n271 m9m10.n270 0.789389
R4329 m9m10.n272 m9m10.n271 0.789389
R4330 m9m10.n273 m9m10.n272 0.789389
R4331 m9m10.n274 m9m10.n273 0.789389
R4332 m9m10.n275 m9m10.n274 0.789389
R4333 m9m10.n276 m9m10.n275 0.789389
R4334 m9m10.n277 m9m10.n276 0.789389
R4335 m9m10.n278 m9m10.n277 0.789389
R4336 m9m10.n279 m9m10.n278 0.789389
R4337 m9m10.n280 m9m10.n279 0.789389
R4338 m9m10.n281 m9m10.n280 0.789389
R4339 m9m10.n282 m9m10.n281 0.789389
R4340 m9m10.n283 m9m10.n282 0.789389
R4341 m9m10.n284 m9m10.n283 0.789389
R4342 m9m10.n285 m9m10.n284 0.789389
R4343 m9m10.n286 m9m10.n285 0.789389
R4344 m9m10.n287 m9m10.n286 0.789389
R4345 m9m10.n288 m9m10.n287 0.789389
R4346 m9m10.n289 m9m10.n288 0.789389
R4347 m9m10.n290 m9m10.n289 0.789389
R4348 m9m10.n291 m9m10.n290 0.789389
R4349 m9m10.n292 m9m10.n291 0.789389
R4350 m9m10.n293 m9m10.n292 0.789389
R4351 m9m10.n294 m9m10.n293 0.789389
R4352 m9m10.n295 m9m10.n294 0.789389
R4353 m9m10.n296 m9m10.n295 0.789389
R4354 m9m10.n297 m9m10.n296 0.789389
R4355 m9m10.n1 m9m10.n0 0.789389
R4356 m9m10.n2 m9m10.n1 0.789389
R4357 m9m10.n3 m9m10.n2 0.789389
R4358 m9m10.n4 m9m10.n3 0.789389
R4359 m9m10.n5 m9m10.n4 0.789389
R4360 m9m10.n6 m9m10.n5 0.789389
R4361 m9m10.n7 m9m10.n6 0.789389
R4362 m9m10.n8 m9m10.n7 0.789389
R4363 m9m10.n9 m9m10.n8 0.789389
R4364 m9m10.n10 m9m10.n9 0.789389
R4365 m9m10.n11 m9m10.n10 0.789389
R4366 m9m10.n12 m9m10.n11 0.789389
R4367 m9m10.n13 m9m10.n12 0.789389
R4368 m9m10.n14 m9m10.n13 0.789389
R4369 m9m10.n15 m9m10.n14 0.789389
R4370 m9m10.n16 m9m10.n15 0.789389
R4371 m9m10.n17 m9m10.n16 0.789389
R4372 m9m10.n18 m9m10.n17 0.789389
R4373 m9m10.n19 m9m10.n18 0.789389
R4374 m9m10.n20 m9m10.n19 0.789389
R4375 m9m10.n21 m9m10.n20 0.789389
R4376 m9m10.n22 m9m10.n21 0.789389
R4377 m9m10.n23 m9m10.n22 0.789389
R4378 m9m10.n24 m9m10.n23 0.789389
R4379 m9m10.n25 m9m10.n24 0.789389
R4380 m9m10.n26 m9m10.n25 0.789389
R4381 m9m10.n27 m9m10.n26 0.789389
R4382 m9m10.n28 m9m10.n27 0.789389
R4383 m9m10.n29 m9m10.n28 0.789389
R4384 m9m10.n30 m9m10.n29 0.789389
R4385 m9m10.n31 m9m10.n30 0.789389
R4386 m9m10.n32 m9m10.n31 0.789389
R4387 m9m10.n33 m9m10.n32 0.789389
R4388 m9m10.n34 m9m10.n33 0.789389
R4389 m9m10.n35 m9m10.n34 0.789389
R4390 m9m10.n36 m9m10.n35 0.789389
R4391 m9m10.n37 m9m10.n36 0.789389
R4392 m9m10.n38 m9m10.n37 0.789389
R4393 m9m10.n39 m9m10.n38 0.789389
R4394 m9m10.n40 m9m10.n39 0.789389
R4395 m9m10.n41 m9m10.n40 0.789389
R4396 m9m10.n42 m9m10.n41 0.789389
R4397 m9m10.n43 m9m10.n42 0.789389
R4398 m9m10.n44 m9m10.n43 0.789389
R4399 m9m10.n45 m9m10.n44 0.789389
R4400 m9m10.n46 m9m10.n45 0.789389
R4401 m9m10.n47 m9m10.n46 0.789389
R4402 m9m10.n48 m9m10.n47 0.789389
R4403 m9m10.n49 m9m10.n48 0.789389
R4404 m9m10.n50 m9m10.n49 0.789389
R4405 m9m10.n51 m9m10.n50 0.789389
R4406 m9m10.n52 m9m10.n51 0.789389
R4407 m9m10.n53 m9m10.n52 0.789389
R4408 m9m10.n54 m9m10.n53 0.789389
R4409 m9m10.n55 m9m10.n54 0.789389
R4410 m9m10.n56 m9m10.n55 0.789389
R4411 m9m10.n57 m9m10.n56 0.789389
R4412 m9m10.n58 m9m10.n57 0.789389
R4413 m9m10.n59 m9m10.n58 0.789389
R4414 m9m10.n60 m9m10.n59 0.789389
R4415 m9m10.n61 m9m10.n60 0.789389
R4416 m9m10.n62 m9m10.n61 0.789389
R4417 m9m10.n63 m9m10.n62 0.789389
R4418 m9m10.n64 m9m10.n63 0.789389
R4419 m9m10.n65 m9m10.n64 0.789389
R4420 m9m10.n66 m9m10.n65 0.789389
R4421 m9m10.n67 m9m10.n66 0.789389
R4422 m9m10.n68 m9m10.n67 0.789389
R4423 m9m10.n69 m9m10.n68 0.789389
R4424 m9m10.n70 m9m10.n69 0.789389
R4425 m9m10.n71 m9m10.n70 0.789389
R4426 m9m10.n72 m9m10.n71 0.789389
R4427 m9m10.n73 m9m10.n72 0.789389
R4428 m9m10.n74 m9m10.n73 0.789389
R4429 m9m10.n75 m9m10.n74 0.789389
R4430 m9m10.n76 m9m10.n75 0.789389
R4431 m9m10.n77 m9m10.n76 0.789389
R4432 m9m10.n78 m9m10.n77 0.789389
R4433 m9m10.n79 m9m10.n78 0.789389
R4434 m9m10.n80 m9m10.n79 0.789389
R4435 m9m10.n81 m9m10.n80 0.789389
R4436 m9m10.n82 m9m10.n81 0.789389
R4437 m9m10.n83 m9m10.n82 0.789389
R4438 m9m10.n84 m9m10.n83 0.789389
R4439 m9m10.n85 m9m10.n84 0.789389
R4440 m9m10.n86 m9m10.n85 0.789389
R4441 m9m10.n87 m9m10.n86 0.789389
R4442 m9m10.n88 m9m10.n87 0.789389
R4443 m9m10.n89 m9m10.n88 0.789389
R4444 m9m10.n90 m9m10.n89 0.789389
R4445 m9m10.n91 m9m10.n90 0.789389
R4446 m9m10.n92 m9m10.n91 0.789389
R4447 m9m10.n93 m9m10.n92 0.789389
R4448 m9m10.n94 m9m10.n93 0.789389
R4449 m9m10.n95 m9m10.n94 0.789389
R4450 m9m10.n96 m9m10.n95 0.789389
R4451 m9m10.n97 m9m10.n96 0.789389
R4452 m9m10.n98 m9m10.n97 0.789389
R4453 m9m10.n197 m9m10.n196 0.789389
R4454 m9m10.n196 m9m10.n195 0.789389
R4455 m9m10.n195 m9m10.n194 0.789389
R4456 m9m10.n194 m9m10.n193 0.789389
R4457 m9m10.n193 m9m10.n192 0.789389
R4458 m9m10.n192 m9m10.n191 0.789389
R4459 m9m10.n191 m9m10.n190 0.789389
R4460 m9m10.n190 m9m10.n189 0.789389
R4461 m9m10.n189 m9m10.n188 0.789389
R4462 m9m10.n188 m9m10.n187 0.789389
R4463 m9m10.n187 m9m10.n186 0.789389
R4464 m9m10.n186 m9m10.n185 0.789389
R4465 m9m10.n185 m9m10.n184 0.789389
R4466 m9m10.n184 m9m10.n183 0.789389
R4467 m9m10.n183 m9m10.n182 0.789389
R4468 m9m10.n182 m9m10.n181 0.789389
R4469 m9m10.n181 m9m10.n180 0.789389
R4470 m9m10.n180 m9m10.n179 0.789389
R4471 m9m10.n179 m9m10.n178 0.789389
R4472 m9m10.n178 m9m10.n177 0.789389
R4473 m9m10.n177 m9m10.n176 0.789389
R4474 m9m10.n176 m9m10.n175 0.789389
R4475 m9m10.n175 m9m10.n174 0.789389
R4476 m9m10.n174 m9m10.n173 0.789389
R4477 m9m10.n173 m9m10.n172 0.789389
R4478 m9m10.n172 m9m10.n171 0.789389
R4479 m9m10.n171 m9m10.n170 0.789389
R4480 m9m10.n170 m9m10.n169 0.789389
R4481 m9m10.n169 m9m10.n168 0.789389
R4482 m9m10.n168 m9m10.n167 0.789389
R4483 m9m10.n167 m9m10.n166 0.789389
R4484 m9m10.n166 m9m10.n165 0.789389
R4485 m9m10.n165 m9m10.n164 0.789389
R4486 m9m10.n164 m9m10.n163 0.789389
R4487 m9m10.n163 m9m10.n162 0.789389
R4488 m9m10.n162 m9m10.n161 0.789389
R4489 m9m10.n161 m9m10.n160 0.789389
R4490 m9m10.n160 m9m10.n159 0.789389
R4491 m9m10.n159 m9m10.n158 0.789389
R4492 m9m10.n158 m9m10.n157 0.789389
R4493 m9m10.n157 m9m10.n156 0.789389
R4494 m9m10.n156 m9m10.n155 0.789389
R4495 m9m10.n155 m9m10.n154 0.789389
R4496 m9m10.n154 m9m10.n153 0.789389
R4497 m9m10.n153 m9m10.n152 0.789389
R4498 m9m10.n152 m9m10.n151 0.789389
R4499 m9m10.n151 m9m10.n150 0.789389
R4500 m9m10.n150 m9m10.n149 0.789389
R4501 m9m10.n149 m9m10.n148 0.789389
R4502 m9m10.n148 m9m10.n147 0.789389
R4503 m9m10.n147 m9m10.n146 0.789389
R4504 m9m10.n146 m9m10.n145 0.789389
R4505 m9m10.n145 m9m10.n144 0.789389
R4506 m9m10.n144 m9m10.n143 0.789389
R4507 m9m10.n143 m9m10.n142 0.789389
R4508 m9m10.n142 m9m10.n141 0.789389
R4509 m9m10.n141 m9m10.n140 0.789389
R4510 m9m10.n140 m9m10.n139 0.789389
R4511 m9m10.n139 m9m10.n138 0.789389
R4512 m9m10.n138 m9m10.n137 0.789389
R4513 m9m10.n137 m9m10.n136 0.789389
R4514 m9m10.n136 m9m10.n135 0.789389
R4515 m9m10.n135 m9m10.n134 0.789389
R4516 m9m10.n134 m9m10.n133 0.789389
R4517 m9m10.n133 m9m10.n132 0.789389
R4518 m9m10.n132 m9m10.n131 0.789389
R4519 m9m10.n131 m9m10.n130 0.789389
R4520 m9m10.n130 m9m10.n129 0.789389
R4521 m9m10.n129 m9m10.n128 0.789389
R4522 m9m10.n128 m9m10.n127 0.789389
R4523 m9m10.n127 m9m10.n126 0.789389
R4524 m9m10.n126 m9m10.n125 0.789389
R4525 m9m10.n125 m9m10.n124 0.789389
R4526 m9m10.n124 m9m10.n123 0.789389
R4527 m9m10.n123 m9m10.n122 0.789389
R4528 m9m10.n122 m9m10.n121 0.789389
R4529 m9m10.n121 m9m10.n120 0.789389
R4530 m9m10.n120 m9m10.n119 0.789389
R4531 m9m10.n119 m9m10.n118 0.789389
R4532 m9m10.n118 m9m10.n117 0.789389
R4533 m9m10.n117 m9m10.n116 0.789389
R4534 m9m10.n116 m9m10.n115 0.789389
R4535 m9m10.n115 m9m10.n114 0.789389
R4536 m9m10.n114 m9m10.n113 0.789389
R4537 m9m10.n113 m9m10.n112 0.789389
R4538 m9m10.n112 m9m10.n111 0.789389
R4539 m9m10.n111 m9m10.n110 0.789389
R4540 m1m2 m1m2.n498 20.1611
R4541 m1m2.n495 m1m2.n494 7.54545
R4542 m1m2.n396 m1m2.t483 6.56346
R4543 m1m2.n297 m1m2.t468 6.56346
R4544 m1m2.n198 m1m2.t162 6.56346
R4545 m1m2.n99 m1m2.t365 6.56346
R4546 m1m2.n0 m1m2.t350 6.56346
R4547 m1m2.n482 m1m2.t116 5.71419
R4548 m1m2.n481 m1m2.t485 5.71419
R4549 m1m2.n480 m1m2.t101 5.71419
R4550 m1m2.n479 m1m2.t229 5.71419
R4551 m1m2.n478 m1m2.t109 5.71419
R4552 m1m2.n477 m1m2.t209 5.71419
R4553 m1m2.n476 m1m2.t472 5.71419
R4554 m1m2.n475 m1m2.t444 5.71419
R4555 m1m2.n474 m1m2.t65 5.71419
R4556 m1m2.n473 m1m2.t309 5.71419
R4557 m1m2.n472 m1m2.t45 5.71419
R4558 m1m2.n471 m1m2.t317 5.71419
R4559 m1m2.n470 m1m2.t54 5.71419
R4560 m1m2.n469 m1m2.t143 5.71419
R4561 m1m2.n468 m1m2.t414 5.71419
R4562 m1m2.n467 m1m2.t390 5.71419
R4563 m1m2.n466 m1m2.t156 5.71419
R4564 m1m2.n465 m1m2.t278 5.71419
R4565 m1m2.n464 m1m2.t489 5.71419
R4566 m1m2.n463 m1m2.t258 5.71419
R4567 m1m2.n462 m1m2.t380 5.71419
R4568 m1m2.n461 m1m2.t266 5.71419
R4569 m1m2.n460 m1m2.t358 5.71419
R4570 m1m2.n459 m1m2.t333 5.71419
R4571 m1m2.n458 m1m2.t96 5.71419
R4572 m1m2.n457 m1m2.t222 5.71419
R4573 m1m2.n456 m1m2.t79 5.71419
R4574 m1m2.n455 m1m2.t204 5.71419
R4575 m1m2.n454 m1m2.t321 5.71419
R4576 m1m2.n453 m1m2.t212 5.71419
R4577 m1m2.n452 m1m2.t301 5.71419
R4578 m1m2.n451 m1m2.t304 5.71419
R4579 m1m2.n450 m1m2.t40 5.71419
R4580 m1m2.n449 m1m2.t161 5.71419
R4581 m1m2.n448 m1m2.t431 5.71419
R4582 m1m2.n447 m1m2.t137 5.71419
R4583 m1m2.n446 m1m2.t409 5.71419
R4584 m1m2.n445 m1m2.t146 5.71419
R4585 m1m2.n444 m1m2.t275 5.71419
R4586 m1m2.n443 m1m2.t245 5.71419
R4587 m1m2.n442 m1m2.t482 5.71419
R4588 m1m2.n441 m1m2.t254 5.71419
R4589 m1m2.n440 m1m2.t374 5.71419
R4590 m1m2.n439 m1m2.t82 5.71419
R4591 m1m2.n438 m1m2.t354 5.71419
R4592 m1m2.n437 m1m2.t470 5.71419
R4593 m1m2.n436 m1m2.t362 5.71419
R4594 m1m2.n435 m1m2.t190 5.71419
R4595 m1m2.n434 m1m2.t427 5.71419
R4596 m1m2.n433 m1m2.t200 5.71419
R4597 m1m2.n432 m1m2.t316 5.71419
R4598 m1m2.n431 m1m2.t180 5.71419
R4599 m1m2.n430 m1m2.t296 5.71419
R4600 m1m2.n429 m1m2.t412 5.71419
R4601 m1m2.n428 m1m2.t305 5.71419
R4602 m1m2.n427 m1m2.t425 5.71419
R4603 m1m2.n426 m1m2.t39 5.71419
R4604 m1m2.n425 m1m2.t284 5.71419
R4605 m1m2.n424 m1m2.t398 5.71419
R4606 m1m2.n423 m1m2.t170 5.71419
R4607 m1m2.n422 m1m2.t386 5.71419
R4608 m1m2.n421 m1m2.t145 5.71419
R4609 m1m2.n420 m1m2.t391 5.71419
R4610 m1m2.n419 m1m2.t3 5.71419
R4611 m1m2.n418 m1m2.t481 5.71419
R4612 m1m2.n417 m1m2.t228 5.71419
R4613 m1m2.n416 m1m2.t491 5.71419
R4614 m1m2.n415 m1m2.t106 5.71419
R4615 m1m2.n414 m1m2.t327 5.71419
R4616 m1m2.n413 m1m2.t89 5.71419
R4617 m1m2.n412 m1m2.t217 5.71419
R4618 m1m2.n411 m1m2.t97 5.71419
R4619 m1m2.n410 m1m2.t447 5.71419
R4620 m1m2.n409 m1m2.t166 5.71419
R4621 m1m2.n408 m1m2.t435 5.71419
R4622 m1m2.n407 m1m2.t51 5.71419
R4623 m1m2.n406 m1m2.t442 5.71419
R4624 m1m2.n405 m1m2.t34 5.71419
R4625 m1m2.n404 m1m2.t150 5.71419
R4626 m1m2.n403 m1m2.t41 5.71419
R4627 m1m2.n402 m1m2.t394 5.71419
R4628 m1m2.n401 m1m2.t131 5.71419
R4629 m1m2.n400 m1m2.t378 5.71419
R4630 m1m2.n399 m1m2.t493 5.71419
R4631 m1m2.n398 m1m2.t263 5.71419
R4632 m1m2.n397 m1m2.t476 5.71419
R4633 m1m2.n396 m1m2.t246 5.71419
R4634 m1m2.n484 m1m2.t497 5.71419
R4635 m1m2.n485 m1m2.t264 5.71419
R4636 m1m2.n486 m1m2.t140 5.71419
R4637 m1m2.n487 m1m2.t285 5.71419
R4638 m1m2.n488 m1m2.t163 5.71419
R4639 m1m2.n489 m1m2.t395 5.71419
R4640 m1m2.n490 m1m2.t153 5.71419
R4641 m1m2.n491 m1m2.t60 5.71419
R4642 m1m2.n492 m1m2.t59 5.71419
R4643 m1m2.n493 m1m2.t323 5.71419
R4644 m1m2.n494 m1m2.t52 5.71419
R4645 m1m2.n513 m1m2.t503 5.71419
R4646 m1m2.n513 m1m2.t524 5.71419
R4647 m1m2.n512 m1m2.t502 5.71419
R4648 m1m2.n512 m1m2.t500 5.71419
R4649 m1m2.n511 m1m2.t528 5.71419
R4650 m1m2.n511 m1m2.t515 5.71419
R4651 m1m2.n510 m1m2.t504 5.71419
R4652 m1m2.n510 m1m2.t523 5.71419
R4653 m1m2.n509 m1m2.t518 5.71419
R4654 m1m2.n509 m1m2.t506 5.71419
R4655 m1m2.n508 m1m2.t510 5.71419
R4656 m1m2.n508 m1m2.t508 5.71419
R4657 m1m2.n507 m1m2.t512 5.71419
R4658 m1m2.n507 m1m2.t501 5.71419
R4659 m1m2.n506 m1m2.t526 5.71419
R4660 m1m2.n506 m1m2.t513 5.71419
R4661 m1m2.n505 m1m2.t514 5.71419
R4662 m1m2.n505 m1m2.t505 5.71419
R4663 m1m2.n504 m1m2.t525 5.71419
R4664 m1m2.n504 m1m2.t516 5.71419
R4665 m1m2.n503 m1m2.t522 5.71419
R4666 m1m2.n503 m1m2.t509 5.71419
R4667 m1m2.n502 m1m2.t519 5.71419
R4668 m1m2.n502 m1m2.t517 5.71419
R4669 m1m2.n501 m1m2.t511 5.71419
R4670 m1m2.n501 m1m2.t529 5.71419
R4671 m1m2.n500 m1m2.t521 5.71419
R4672 m1m2.n500 m1m2.t520 5.71419
R4673 m1m2.n499 m1m2.t507 5.71419
R4674 m1m2.n499 m1m2.t527 5.71419
R4675 m1m2.n395 m1m2.t92 5.71419
R4676 m1m2.n394 m1m2.t369 5.71419
R4677 m1m2.n393 m1m2.t100 5.71419
R4678 m1m2.n392 m1m2.t102 5.71419
R4679 m1m2.n391 m1m2.t203 5.71419
R4680 m1m2.n390 m1m2.t438 5.71419
R4681 m1m2.n389 m1m2.t211 5.71419
R4682 m1m2.n388 m1m2.t328 5.71419
R4683 m1m2.n387 m1m2.t192 5.71419
R4684 m1m2.n386 m1m2.t308 5.71419
R4685 m1m2.n385 m1m2.t44 5.71419
R4686 m1m2.n384 m1m2.t46 5.71419
R4687 m1m2.n383 m1m2.t169 5.71419
R4688 m1m2.n382 m1m2.t28 5.71419
R4689 m1m2.n381 m1m2.t144 5.71419
R4690 m1m2.n380 m1m2.t271 5.71419
R4691 m1m2.n379 m1m2.t155 5.71419
R4692 m1m2.n378 m1m2.t249 5.71419
R4693 m1m2.n377 m1m2.t12 5.71419
R4694 m1m2.n376 m1m2.t490 5.71419
R4695 m1m2.n375 m1m2.t105 5.71419
R4696 m1m2.n374 m1m2.t351 5.71419
R4697 m1m2.n373 m1m2.t88 5.71419
R4698 m1m2.n372 m1m2.t360 5.71419
R4699 m1m2.n371 m1m2.t95 5.71419
R4700 m1m2.n370 m1m2.t196 5.71419
R4701 m1m2.n369 m1m2.t456 5.71419
R4702 m1m2.n368 m1m2.t434 5.71419
R4703 m1m2.n367 m1m2.t205 5.71419
R4704 m1m2.n366 m1m2.t322 5.71419
R4705 m1m2.n365 m1m2.t33 5.71419
R4706 m1m2.n364 m1m2.t303 5.71419
R4707 m1m2.n363 m1m2.t421 5.71419
R4708 m1m2.n362 m1m2.t311 5.71419
R4709 m1m2.n361 m1m2.t401 5.71419
R4710 m1m2.n360 m1m2.t377 5.71419
R4711 m1m2.n359 m1m2.t138 5.71419
R4712 m1m2.n358 m1m2.t262 5.71419
R4713 m1m2.n357 m1m2.t120 5.71419
R4714 m1m2.n356 m1m2.t244 5.71419
R4715 m1m2.n355 m1m2.t367 5.71419
R4716 m1m2.n354 m1m2.t253 5.71419
R4717 m1m2.n353 m1m2.t342 5.71419
R4718 m1m2.n352 m1m2.t343 5.71419
R4719 m1m2.n351 m1m2.t83 5.71419
R4720 m1m2.n350 m1m2.t208 5.71419
R4721 m1m2.n349 m1m2.t471 5.71419
R4722 m1m2.n348 m1m2.t189 5.71419
R4723 m1m2.n347 m1m2.t449 5.71419
R4724 m1m2.n346 m1m2.t199 5.71419
R4725 m1m2.n345 m1m2.t314 5.71419
R4726 m1m2.n344 m1m2.t290 5.71419
R4727 m1m2.n343 m1m2.t24 5.71419
R4728 m1m2.n342 m1m2.t297 5.71419
R4729 m1m2.n341 m1m2.t413 5.71419
R4730 m1m2.n340 m1m2.t126 5.71419
R4731 m1m2.n339 m1m2.t397 5.71419
R4732 m1m2.n338 m1m2.t9 5.71419
R4733 m1m2.n337 m1m2.t403 5.71419
R4734 m1m2.n336 m1m2.t235 5.71419
R4735 m1m2.n335 m1m2.t467 5.71419
R4736 m1m2.n334 m1m2.t241 5.71419
R4737 m1m2.n333 m1m2.t357 5.71419
R4738 m1m2.n332 m1m2.t225 5.71419
R4739 m1m2.n331 m1m2.t338 5.71419
R4740 m1m2.n330 m1m2.t453 5.71419
R4741 m1m2.n329 m1m2.t346 5.71419
R4742 m1m2.n328 m1m2.t462 5.71419
R4743 m1m2.n327 m1m2.t23 5.71419
R4744 m1m2.n326 m1m2.t270 5.71419
R4745 m1m2.n325 m1m2.t388 5.71419
R4746 m1m2.n324 m1m2.t152 5.71419
R4747 m1m2.n323 m1m2.t372 5.71419
R4748 m1m2.n322 m1m2.t130 5.71419
R4749 m1m2.n321 m1m2.t379 5.71419
R4750 m1m2.n320 m1m2.t494 5.71419
R4751 m1m2.n319 m1m2.t466 5.71419
R4752 m1m2.n318 m1m2.t215 5.71419
R4753 m1m2.n317 m1m2.t478 5.71419
R4754 m1m2.n316 m1m2.t93 5.71419
R4755 m1m2.n315 m1m2.t312 5.71419
R4756 m1m2.n314 m1m2.t76 5.71419
R4757 m1m2.n313 m1m2.t202 5.71419
R4758 m1m2.n312 m1m2.t85 5.71419
R4759 m1m2.n311 m1m2.t439 5.71419
R4760 m1m2.n310 m1m2.t149 5.71419
R4761 m1m2.n309 m1m2.t420 5.71419
R4762 m1m2.n308 m1m2.t37 5.71419
R4763 m1m2.n307 m1m2.t430 5.71419
R4764 m1m2.n306 m1m2.t17 5.71419
R4765 m1m2.n305 m1m2.t135 5.71419
R4766 m1m2.n304 m1m2.t25 5.71419
R4767 m1m2.n303 m1m2.t385 5.71419
R4768 m1m2.n302 m1m2.t118 5.71419
R4769 m1m2.n301 m1m2.t366 5.71419
R4770 m1m2.n300 m1m2.t480 5.71419
R4771 m1m2.n299 m1m2.t250 5.71419
R4772 m1m2.n298 m1m2.t459 5.71419
R4773 m1m2.n297 m1m2.t236 5.71419
R4774 m1m2.n296 m1m2.t428 5.71419
R4775 m1m2.n295 m1m2.t201 5.71419
R4776 m1m2.n294 m1m2.t436 5.71419
R4777 m1m2.n293 m1m2.t437 5.71419
R4778 m1m2.n292 m1m2.t26 5.71419
R4779 m1m2.n291 m1m2.t273 5.71419
R4780 m1m2.n290 m1m2.t36 5.71419
R4781 m1m2.n289 m1m2.t154 5.71419
R4782 m1m2.n288 m1m2.t14 5.71419
R4783 m1m2.n287 m1m2.t132 5.71419
R4784 m1m2.n286 m1m2.t381 5.71419
R4785 m1m2.n285 m1m2.t382 5.71419
R4786 m1m2.n284 m1m2.t495 5.71419
R4787 m1m2.n283 m1m2.t361 5.71419
R4788 m1m2.n282 m1m2.t479 5.71419
R4789 m1m2.n281 m1m2.t94 5.71419
R4790 m1m2.n280 m1m2.t486 5.71419
R4791 m1m2.n279 m1m2.t77 5.71419
R4792 m1m2.n278 m1m2.t348 5.71419
R4793 m1m2.n277 m1m2.t324 5.71419
R4794 m1m2.n276 m1m2.t440 5.71419
R4795 m1m2.n275 m1m2.t186 5.71419
R4796 m1m2.n274 m1m2.t422 5.71419
R4797 m1m2.n273 m1m2.t195 5.71419
R4798 m1m2.n272 m1m2.t432 5.71419
R4799 m1m2.n271 m1m2.t18 5.71419
R4800 m1m2.n270 m1m2.t293 5.71419
R4801 m1m2.n269 m1m2.t265 5.71419
R4802 m1m2.n268 m1m2.t30 5.71419
R4803 m1m2.n267 m1m2.t147 5.71419
R4804 m1m2.n266 m1m2.t368 5.71419
R4805 m1m2.n265 m1m2.t129 5.71419
R4806 m1m2.n264 m1m2.t252 5.71419
R4807 m1m2.n263 m1m2.t134 5.71419
R4808 m1m2.n262 m1m2.t237 5.71419
R4809 m1m2.n261 m1m2.t210 5.71419
R4810 m1m2.n260 m1m2.t473 5.71419
R4811 m1m2.n259 m1m2.t90 5.71419
R4812 m1m2.n258 m1m2.t450 5.71419
R4813 m1m2.n257 m1m2.t73 5.71419
R4814 m1m2.n256 m1m2.t198 5.71419
R4815 m1m2.n255 m1m2.t80 5.71419
R4816 m1m2.n254 m1m2.t178 5.71419
R4817 m1m2.n253 m1m2.t181 5.71419
R4818 m1m2.n252 m1m2.t415 5.71419
R4819 m1m2.n251 m1m2.t35 5.71419
R4820 m1m2.n250 m1m2.t306 5.71419
R4821 m1m2.n249 m1m2.t11 5.71419
R4822 m1m2.n248 m1m2.t288 5.71419
R4823 m1m2.n247 m1m2.t21 5.71419
R4824 m1m2.n246 m1m2.t141 5.71419
R4825 m1m2.n245 m1m2.t114 5.71419
R4826 m1m2.n244 m1m2.t359 5.71419
R4827 m1m2.n243 m1m2.t122 5.71419
R4828 m1m2.n242 m1m2.t247 5.71419
R4829 m1m2.n241 m1m2.t455 5.71419
R4830 m1m2.n240 m1m2.t233 5.71419
R4831 m1m2.n239 m1m2.t345 5.71419
R4832 m1m2.n238 m1m2.t239 5.71419
R4833 m1m2.n237 m1m2.t62 5.71419
R4834 m1m2.n236 m1m2.t302 5.71419
R4835 m1m2.n235 m1m2.t70 5.71419
R4836 m1m2.n234 m1m2.t193 5.71419
R4837 m1m2.n233 m1m2.t50 5.71419
R4838 m1m2.n232 m1m2.t174 5.71419
R4839 m1m2.n231 m1m2.t292 5.71419
R4840 m1m2.n230 m1m2.t183 5.71419
R4841 m1m2.n229 m1m2.t298 5.71419
R4842 m1m2.n228 m1m2.t221 5.71419
R4843 m1m2.n227 m1m2.t451 5.71419
R4844 m1m2.n226 m1m2.t74 5.71419
R4845 m1m2.n225 m1m2.t341 5.71419
R4846 m1m2.n224 m1m2.t58 5.71419
R4847 m1m2.n223 m1m2.t329 5.71419
R4848 m1m2.n222 m1m2.t66 5.71419
R4849 m1m2.n221 m1m2.t188 5.71419
R4850 m1m2.n220 m1m2.t160 5.71419
R4851 m1m2.n219 m1m2.t399 5.71419
R4852 m1m2.n218 m1m2.t171 5.71419
R4853 m1m2.n217 m1m2.t289 5.71419
R4854 m1m2.n216 m1m2.t496 5.71419
R4855 m1m2.n215 m1m2.t274 5.71419
R4856 m1m2.n214 m1m2.t389 5.71419
R4857 m1m2.n213 m1m2.t279 5.71419
R4858 m1m2.n212 m1m2.t124 5.71419
R4859 m1m2.n211 m1m2.t339 5.71419
R4860 m1m2.n210 m1m2.t107 5.71419
R4861 m1m2.n209 m1m2.t234 5.71419
R4862 m1m2.n208 m1m2.t113 5.71419
R4863 m1m2.n207 m1m2.t218 5.71419
R4864 m1m2.n206 m1m2.t332 5.71419
R4865 m1m2.n205 m1m2.t223 5.71419
R4866 m1m2.n204 m1m2.t72 5.71419
R4867 m1m2.n203 m1m2.t315 5.71419
R4868 m1m2.n202 m1m2.t53 5.71419
R4869 m1m2.n201 m1m2.t176 5.71419
R4870 m1m2.n200 m1m2.t441 5.71419
R4871 m1m2.n199 m1m2.t151 5.71419
R4872 m1m2.n198 m1m2.t424 5.71419
R4873 m1m2.n197 m1m2.t411 5.71419
R4874 m1m2.n196 m1m2.t187 5.71419
R4875 m1m2.n195 m1m2.t423 5.71419
R4876 m1m2.n194 m1m2.t426 5.71419
R4877 m1m2.n193 m1m2.t10 5.71419
R4878 m1m2.n192 m1m2.t257 5.71419
R4879 m1m2.n191 m1m2.t20 5.71419
R4880 m1m2.n190 m1m2.t139 5.71419
R4881 m1m2.n189 m1m2.t2 5.71419
R4882 m1m2.n188 m1m2.t121 5.71419
R4883 m1m2.n187 m1m2.t370 5.71419
R4884 m1m2.n186 m1m2.t371 5.71419
R4885 m1m2.n185 m1m2.t484 5.71419
R4886 m1m2.n184 m1m2.t347 5.71419
R4887 m1m2.n183 m1m2.t463 5.71419
R4888 m1m2.n182 m1m2.t84 5.71419
R4889 m1m2.n181 m1m2.t474 5.71419
R4890 m1m2.n180 m1m2.t68 5.71419
R4891 m1m2.n179 m1m2.t337 5.71419
R4892 m1m2.n178 m1m2.t310 5.71419
R4893 m1m2.n177 m1m2.t429 5.71419
R4894 m1m2.n176 m1m2.t173 5.71419
R4895 m1m2.n175 m1m2.t407 5.71419
R4896 m1m2.n174 m1m2.t182 5.71419
R4897 m1m2.n173 m1m2.t416 5.71419
R4898 m1m2.n172 m1m2.t4 5.71419
R4899 m1m2.n171 m1m2.t283 5.71419
R4900 m1m2.n170 m1m2.t251 5.71419
R4901 m1m2.n169 m1m2.t15 5.71419
R4902 m1m2.n168 m1m2.t133 5.71419
R4903 m1m2.n167 m1m2.t352 5.71419
R4904 m1m2.n166 m1m2.t115 5.71419
R4905 m1m2.n165 m1m2.t242 5.71419
R4906 m1m2.n164 m1m2.t123 5.71419
R4907 m1m2.n163 m1m2.t226 5.71419
R4908 m1m2.n162 m1m2.t197 5.71419
R4909 m1m2.n161 m1m2.t458 5.71419
R4910 m1m2.n160 m1m2.t78 5.71419
R4911 m1m2.n159 m1m2.t443 5.71419
R4912 m1m2.n158 m1m2.t63 5.71419
R4913 m1m2.n157 m1m2.t184 5.71419
R4914 m1m2.n156 m1m2.t71 5.71419
R4915 m1m2.n155 m1m2.t164 5.71419
R4916 m1m2.n154 m1m2.t167 5.71419
R4917 m1m2.n153 m1m2.t402 5.71419
R4918 m1m2.n152 m1m2.t19 5.71419
R4919 m1m2.n151 m1m2.t294 5.71419
R4920 m1m2.n150 m1m2.t0 5.71419
R4921 m1m2.n149 m1m2.t277 5.71419
R4922 m1m2.n148 m1m2.t6 5.71419
R4923 m1m2.n147 m1m2.t128 5.71419
R4924 m1m2.n146 m1m2.t104 5.71419
R4925 m1m2.n145 m1m2.t344 5.71419
R4926 m1m2.n144 m1m2.t112 5.71419
R4927 m1m2.n143 m1m2.t238 5.71419
R4928 m1m2.n142 m1m2.t445 5.71419
R4929 m1m2.n141 m1m2.t220 5.71419
R4930 m1m2.n140 m1m2.t335 5.71419
R4931 m1m2.n139 m1m2.t230 5.71419
R4932 m1m2.n138 m1m2.t48 5.71419
R4933 m1m2.n137 m1m2.t291 5.71419
R4934 m1m2.n136 m1m2.t57 5.71419
R4935 m1m2.n135 m1m2.t179 5.71419
R4936 m1m2.n134 m1m2.t38 5.71419
R4937 m1m2.n133 m1m2.t158 5.71419
R4938 m1m2.n132 m1m2.t281 5.71419
R4939 m1m2.n131 m1m2.t168 5.71419
R4940 m1m2.n130 m1m2.t287 5.71419
R4941 m1m2.n129 m1m2.t418 5.71419
R4942 m1m2.n128 m1m2.t157 5.71419
R4943 m1m2.n127 m1m2.t280 5.71419
R4944 m1m2.n126 m1m2.t43 5.71419
R4945 m1m2.n125 m1m2.t260 5.71419
R4946 m1m2.n124 m1m2.t22 5.71419
R4947 m1m2.n123 m1m2.t269 5.71419
R4948 m1m2.n122 m1m2.t387 5.71419
R4949 m1m2.n121 m1m2.t364 5.71419
R4950 m1m2.n120 m1m2.t98 5.71419
R4951 m1m2.n119 m1m2.t373 5.71419
R4952 m1m2.n118 m1m2.t487 5.71419
R4953 m1m2.n117 m1m2.t206 5.71419
R4954 m1m2.n116 m1m2.t465 5.71419
R4955 m1m2.n115 m1m2.t87 5.71419
R4956 m1m2.n114 m1m2.t477 5.71419
R4957 m1m2.n113 m1m2.t330 5.71419
R4958 m1m2.n112 m1m2.t42 5.71419
R4959 m1m2.n111 m1m2.t313 5.71419
R4960 m1m2.n110 m1m2.t433 5.71419
R4961 m1m2.n109 m1m2.t320 5.71419
R4962 m1m2.n108 m1m2.t410 5.71419
R4963 m1m2.n107 m1m2.t31 5.71419
R4964 m1m2.n106 m1m2.t419 5.71419
R4965 m1m2.n105 m1m2.t276 5.71419
R4966 m1m2.n104 m1m2.t7 5.71419
R4967 m1m2.n103 m1m2.t255 5.71419
R4968 m1m2.n102 m1m2.t375 5.71419
R4969 m1m2.n101 m1m2.t136 5.71419
R4970 m1m2.n100 m1m2.t355 5.71419
R4971 m1m2.n99 m1m2.t117 5.71419
R4972 m1m2.n98 m1m2.t454 5.71419
R4973 m1m2.n97 m1m2.t232 5.71419
R4974 m1m2.n96 m1m2.t461 5.71419
R4975 m1m2.n95 m1m2.t464 5.71419
R4976 m1m2.n94 m1m2.t61 5.71419
R4977 m1m2.n93 m1m2.t300 5.71419
R4978 m1m2.n92 m1m2.t69 5.71419
R4979 m1m2.n91 m1m2.t191 5.71419
R4980 m1m2.n90 m1m2.t49 5.71419
R4981 m1m2.n89 m1m2.t172 5.71419
R4982 m1m2.n88 m1m2.t406 5.71419
R4983 m1m2.n87 m1m2.t408 5.71419
R4984 m1m2.n86 m1m2.t27 5.71419
R4985 m1m2.n85 m1m2.t393 5.71419
R4986 m1m2.n84 m1m2.t5 5.71419
R4987 m1m2.n83 m1m2.t127 5.71419
R4988 m1m2.n82 m1m2.t13 5.71419
R4989 m1m2.n81 m1m2.t110 5.71419
R4990 m1m2.n80 m1m2.t384 5.71419
R4991 m1m2.n79 m1m2.t353 5.71419
R4992 m1m2.n78 m1m2.t469 5.71419
R4993 m1m2.n77 m1m2.t219 5.71419
R4994 m1m2.n76 m1m2.t448 5.71419
R4995 m1m2.n75 m1m2.t227 5.71419
R4996 m1m2.n74 m1m2.t457 5.71419
R4997 m1m2.n73 m1m2.t55 5.71419
R4998 m1m2.n72 m1m2.t326 5.71419
R4999 m1m2.n71 m1m2.t295 5.71419
R5000 m1m2.n70 m1m2.t64 5.71419
R5001 m1m2.n69 m1m2.t185 5.71419
R5002 m1m2.n68 m1m2.t396 5.71419
R5003 m1m2.n67 m1m2.t165 5.71419
R5004 m1m2.n66 m1m2.t286 5.71419
R5005 m1m2.n65 m1m2.t175 5.71419
R5006 m1m2.n64 m1m2.t268 5.71419
R5007 m1m2.n63 m1m2.t240 5.71419
R5008 m1m2.n62 m1m2.t1 5.71419
R5009 m1m2.n61 m1m2.t119 5.71419
R5010 m1m2.n60 m1m2.t488 5.71419
R5011 m1m2.n59 m1m2.t103 5.71419
R5012 m1m2.n58 m1m2.t231 5.71419
R5013 m1m2.n57 m1m2.t111 5.71419
R5014 m1m2.n56 m1m2.t213 5.71419
R5015 m1m2.n55 m1m2.t214 5.71419
R5016 m1m2.n54 m1m2.t446 5.71419
R5017 m1m2.n53 m1m2.t67 5.71419
R5018 m1m2.n52 m1m2.t336 5.71419
R5019 m1m2.n51 m1m2.t47 5.71419
R5020 m1m2.n50 m1m2.t319 5.71419
R5021 m1m2.n49 m1m2.t56 5.71419
R5022 m1m2.n48 m1m2.t177 5.71419
R5023 m1m2.n47 m1m2.t148 5.71419
R5024 m1m2.n46 m1m2.t392 5.71419
R5025 m1m2.n45 m1m2.t159 5.71419
R5026 m1m2.n44 m1m2.t282 5.71419
R5027 m1m2.n43 m1m2.t492 5.71419
R5028 m1m2.n42 m1m2.t261 5.71419
R5029 m1m2.n41 m1m2.t383 5.71419
R5030 m1m2.n40 m1m2.t272 5.71419
R5031 m1m2.n39 m1m2.t91 5.71419
R5032 m1m2.n38 m1m2.t334 5.71419
R5033 m1m2.n37 m1m2.t99 5.71419
R5034 m1m2.n36 m1m2.t224 5.71419
R5035 m1m2.n35 m1m2.t81 5.71419
R5036 m1m2.n34 m1m2.t207 5.71419
R5037 m1m2.n33 m1m2.t325 5.71419
R5038 m1m2.n32 m1m2.t216 5.71419
R5039 m1m2.n31 m1m2.t331 5.71419
R5040 m1m2.n30 m1m2.t404 5.71419
R5041 m1m2.n29 m1m2.t142 5.71419
R5042 m1m2.n28 m1m2.t267 5.71419
R5043 m1m2.n27 m1m2.t32 5.71419
R5044 m1m2.n26 m1m2.t248 5.71419
R5045 m1m2.n25 m1m2.t8 5.71419
R5046 m1m2.n24 m1m2.t256 5.71419
R5047 m1m2.n23 m1m2.t376 5.71419
R5048 m1m2.n22 m1m2.t349 5.71419
R5049 m1m2.n21 m1m2.t86 5.71419
R5050 m1m2.n20 m1m2.t356 5.71419
R5051 m1m2.n19 m1m2.t475 5.71419
R5052 m1m2.n18 m1m2.t194 5.71419
R5053 m1m2.n17 m1m2.t452 5.71419
R5054 m1m2.n16 m1m2.t75 5.71419
R5055 m1m2.n15 m1m2.t460 5.71419
R5056 m1m2.n14 m1m2.t318 5.71419
R5057 m1m2.n13 m1m2.t29 5.71419
R5058 m1m2.n12 m1m2.t299 5.71419
R5059 m1m2.n11 m1m2.t417 5.71419
R5060 m1m2.n10 m1m2.t307 5.71419
R5061 m1m2.n9 m1m2.t400 5.71419
R5062 m1m2.n8 m1m2.t16 5.71419
R5063 m1m2.n7 m1m2.t405 5.71419
R5064 m1m2.n6 m1m2.t259 5.71419
R5065 m1m2.n5 m1m2.t498 5.71419
R5066 m1m2.n4 m1m2.t243 5.71419
R5067 m1m2.n3 m1m2.t363 5.71419
R5068 m1m2.n2 m1m2.t125 5.71419
R5069 m1m2.n1 m1m2.t340 5.71419
R5070 m1m2.n0 m1m2.t108 5.71419
R5071 m1m2.n483 m1m2.t499 5.71419
R5072 m1m2.n496 m1m2.n495 4.5005
R5073 m1m2.n497 m1m2.n496 4.5005
R5074 m1m2.n498 m1m2.n497 4.5005
R5075 m1m2 m1m2.n513 4.03574
R5076 m1m2.n495 m1m2.n395 3.04545
R5077 m1m2.n496 m1m2.n296 3.04545
R5078 m1m2.n497 m1m2.n197 3.04545
R5079 m1m2.n498 m1m2.n98 2.98587
R5080 m1m2.n397 m1m2.n396 0.849769
R5081 m1m2.n398 m1m2.n397 0.849769
R5082 m1m2.n399 m1m2.n398 0.849769
R5083 m1m2.n400 m1m2.n399 0.849769
R5084 m1m2.n401 m1m2.n400 0.849769
R5085 m1m2.n402 m1m2.n401 0.849769
R5086 m1m2.n403 m1m2.n402 0.849769
R5087 m1m2.n404 m1m2.n403 0.849769
R5088 m1m2.n405 m1m2.n404 0.849769
R5089 m1m2.n406 m1m2.n405 0.849769
R5090 m1m2.n407 m1m2.n406 0.849769
R5091 m1m2.n408 m1m2.n407 0.849769
R5092 m1m2.n409 m1m2.n408 0.849769
R5093 m1m2.n410 m1m2.n409 0.849769
R5094 m1m2.n411 m1m2.n410 0.849769
R5095 m1m2.n412 m1m2.n411 0.849769
R5096 m1m2.n413 m1m2.n412 0.849769
R5097 m1m2.n414 m1m2.n413 0.849769
R5098 m1m2.n415 m1m2.n414 0.849769
R5099 m1m2.n416 m1m2.n415 0.849769
R5100 m1m2.n417 m1m2.n416 0.849769
R5101 m1m2.n418 m1m2.n417 0.849769
R5102 m1m2.n419 m1m2.n418 0.849769
R5103 m1m2.n420 m1m2.n419 0.849769
R5104 m1m2.n421 m1m2.n420 0.849769
R5105 m1m2.n422 m1m2.n421 0.849769
R5106 m1m2.n423 m1m2.n422 0.849769
R5107 m1m2.n424 m1m2.n423 0.849769
R5108 m1m2.n425 m1m2.n424 0.849769
R5109 m1m2.n426 m1m2.n425 0.849769
R5110 m1m2.n427 m1m2.n426 0.849769
R5111 m1m2.n428 m1m2.n427 0.849769
R5112 m1m2.n429 m1m2.n428 0.849769
R5113 m1m2.n430 m1m2.n429 0.849769
R5114 m1m2.n431 m1m2.n430 0.849769
R5115 m1m2.n432 m1m2.n431 0.849769
R5116 m1m2.n433 m1m2.n432 0.849769
R5117 m1m2.n434 m1m2.n433 0.849769
R5118 m1m2.n435 m1m2.n434 0.849769
R5119 m1m2.n436 m1m2.n435 0.849769
R5120 m1m2.n437 m1m2.n436 0.849769
R5121 m1m2.n438 m1m2.n437 0.849769
R5122 m1m2.n439 m1m2.n438 0.849769
R5123 m1m2.n440 m1m2.n439 0.849769
R5124 m1m2.n441 m1m2.n440 0.849769
R5125 m1m2.n442 m1m2.n441 0.849769
R5126 m1m2.n443 m1m2.n442 0.849769
R5127 m1m2.n444 m1m2.n443 0.849769
R5128 m1m2.n445 m1m2.n444 0.849769
R5129 m1m2.n446 m1m2.n445 0.849769
R5130 m1m2.n447 m1m2.n446 0.849769
R5131 m1m2.n448 m1m2.n447 0.849769
R5132 m1m2.n449 m1m2.n448 0.849769
R5133 m1m2.n450 m1m2.n449 0.849769
R5134 m1m2.n451 m1m2.n450 0.849769
R5135 m1m2.n452 m1m2.n451 0.849769
R5136 m1m2.n453 m1m2.n452 0.849769
R5137 m1m2.n454 m1m2.n453 0.849769
R5138 m1m2.n455 m1m2.n454 0.849769
R5139 m1m2.n456 m1m2.n455 0.849769
R5140 m1m2.n457 m1m2.n456 0.849769
R5141 m1m2.n458 m1m2.n457 0.849769
R5142 m1m2.n459 m1m2.n458 0.849769
R5143 m1m2.n460 m1m2.n459 0.849769
R5144 m1m2.n461 m1m2.n460 0.849769
R5145 m1m2.n462 m1m2.n461 0.849769
R5146 m1m2.n463 m1m2.n462 0.849769
R5147 m1m2.n464 m1m2.n463 0.849769
R5148 m1m2.n465 m1m2.n464 0.849769
R5149 m1m2.n466 m1m2.n465 0.849769
R5150 m1m2.n467 m1m2.n466 0.849769
R5151 m1m2.n468 m1m2.n467 0.849769
R5152 m1m2.n469 m1m2.n468 0.849769
R5153 m1m2.n470 m1m2.n469 0.849769
R5154 m1m2.n471 m1m2.n470 0.849769
R5155 m1m2.n472 m1m2.n471 0.849769
R5156 m1m2.n473 m1m2.n472 0.849769
R5157 m1m2.n474 m1m2.n473 0.849769
R5158 m1m2.n475 m1m2.n474 0.849769
R5159 m1m2.n476 m1m2.n475 0.849769
R5160 m1m2.n477 m1m2.n476 0.849769
R5161 m1m2.n478 m1m2.n477 0.849769
R5162 m1m2.n479 m1m2.n478 0.849769
R5163 m1m2.n480 m1m2.n479 0.849769
R5164 m1m2.n481 m1m2.n480 0.849769
R5165 m1m2.n482 m1m2.n481 0.849769
R5166 m1m2.n483 m1m2.n482 0.849769
R5167 m1m2.n298 m1m2.n297 0.849769
R5168 m1m2.n299 m1m2.n298 0.849769
R5169 m1m2.n300 m1m2.n299 0.849769
R5170 m1m2.n301 m1m2.n300 0.849769
R5171 m1m2.n302 m1m2.n301 0.849769
R5172 m1m2.n303 m1m2.n302 0.849769
R5173 m1m2.n304 m1m2.n303 0.849769
R5174 m1m2.n305 m1m2.n304 0.849769
R5175 m1m2.n306 m1m2.n305 0.849769
R5176 m1m2.n307 m1m2.n306 0.849769
R5177 m1m2.n308 m1m2.n307 0.849769
R5178 m1m2.n309 m1m2.n308 0.849769
R5179 m1m2.n310 m1m2.n309 0.849769
R5180 m1m2.n311 m1m2.n310 0.849769
R5181 m1m2.n312 m1m2.n311 0.849769
R5182 m1m2.n313 m1m2.n312 0.849769
R5183 m1m2.n314 m1m2.n313 0.849769
R5184 m1m2.n315 m1m2.n314 0.849769
R5185 m1m2.n316 m1m2.n315 0.849769
R5186 m1m2.n317 m1m2.n316 0.849769
R5187 m1m2.n318 m1m2.n317 0.849769
R5188 m1m2.n319 m1m2.n318 0.849769
R5189 m1m2.n320 m1m2.n319 0.849769
R5190 m1m2.n321 m1m2.n320 0.849769
R5191 m1m2.n322 m1m2.n321 0.849769
R5192 m1m2.n323 m1m2.n322 0.849769
R5193 m1m2.n324 m1m2.n323 0.849769
R5194 m1m2.n325 m1m2.n324 0.849769
R5195 m1m2.n326 m1m2.n325 0.849769
R5196 m1m2.n327 m1m2.n326 0.849769
R5197 m1m2.n328 m1m2.n327 0.849769
R5198 m1m2.n329 m1m2.n328 0.849769
R5199 m1m2.n330 m1m2.n329 0.849769
R5200 m1m2.n331 m1m2.n330 0.849769
R5201 m1m2.n332 m1m2.n331 0.849769
R5202 m1m2.n333 m1m2.n332 0.849769
R5203 m1m2.n334 m1m2.n333 0.849769
R5204 m1m2.n335 m1m2.n334 0.849769
R5205 m1m2.n336 m1m2.n335 0.849769
R5206 m1m2.n337 m1m2.n336 0.849769
R5207 m1m2.n338 m1m2.n337 0.849769
R5208 m1m2.n339 m1m2.n338 0.849769
R5209 m1m2.n340 m1m2.n339 0.849769
R5210 m1m2.n341 m1m2.n340 0.849769
R5211 m1m2.n342 m1m2.n341 0.849769
R5212 m1m2.n343 m1m2.n342 0.849769
R5213 m1m2.n344 m1m2.n343 0.849769
R5214 m1m2.n345 m1m2.n344 0.849769
R5215 m1m2.n346 m1m2.n345 0.849769
R5216 m1m2.n347 m1m2.n346 0.849769
R5217 m1m2.n348 m1m2.n347 0.849769
R5218 m1m2.n349 m1m2.n348 0.849769
R5219 m1m2.n350 m1m2.n349 0.849769
R5220 m1m2.n351 m1m2.n350 0.849769
R5221 m1m2.n352 m1m2.n351 0.849769
R5222 m1m2.n353 m1m2.n352 0.849769
R5223 m1m2.n354 m1m2.n353 0.849769
R5224 m1m2.n355 m1m2.n354 0.849769
R5225 m1m2.n356 m1m2.n355 0.849769
R5226 m1m2.n357 m1m2.n356 0.849769
R5227 m1m2.n358 m1m2.n357 0.849769
R5228 m1m2.n359 m1m2.n358 0.849769
R5229 m1m2.n360 m1m2.n359 0.849769
R5230 m1m2.n361 m1m2.n360 0.849769
R5231 m1m2.n362 m1m2.n361 0.849769
R5232 m1m2.n363 m1m2.n362 0.849769
R5233 m1m2.n364 m1m2.n363 0.849769
R5234 m1m2.n365 m1m2.n364 0.849769
R5235 m1m2.n366 m1m2.n365 0.849769
R5236 m1m2.n367 m1m2.n366 0.849769
R5237 m1m2.n368 m1m2.n367 0.849769
R5238 m1m2.n369 m1m2.n368 0.849769
R5239 m1m2.n370 m1m2.n369 0.849769
R5240 m1m2.n371 m1m2.n370 0.849769
R5241 m1m2.n372 m1m2.n371 0.849769
R5242 m1m2.n373 m1m2.n372 0.849769
R5243 m1m2.n374 m1m2.n373 0.849769
R5244 m1m2.n375 m1m2.n374 0.849769
R5245 m1m2.n376 m1m2.n375 0.849769
R5246 m1m2.n377 m1m2.n376 0.849769
R5247 m1m2.n378 m1m2.n377 0.849769
R5248 m1m2.n379 m1m2.n378 0.849769
R5249 m1m2.n380 m1m2.n379 0.849769
R5250 m1m2.n381 m1m2.n380 0.849769
R5251 m1m2.n382 m1m2.n381 0.849769
R5252 m1m2.n383 m1m2.n382 0.849769
R5253 m1m2.n384 m1m2.n383 0.849769
R5254 m1m2.n385 m1m2.n384 0.849769
R5255 m1m2.n386 m1m2.n385 0.849769
R5256 m1m2.n387 m1m2.n386 0.849769
R5257 m1m2.n388 m1m2.n387 0.849769
R5258 m1m2.n389 m1m2.n388 0.849769
R5259 m1m2.n390 m1m2.n389 0.849769
R5260 m1m2.n391 m1m2.n390 0.849769
R5261 m1m2.n392 m1m2.n391 0.849769
R5262 m1m2.n393 m1m2.n392 0.849769
R5263 m1m2.n394 m1m2.n393 0.849769
R5264 m1m2.n395 m1m2.n394 0.849769
R5265 m1m2.n199 m1m2.n198 0.849769
R5266 m1m2.n200 m1m2.n199 0.849769
R5267 m1m2.n201 m1m2.n200 0.849769
R5268 m1m2.n202 m1m2.n201 0.849769
R5269 m1m2.n203 m1m2.n202 0.849769
R5270 m1m2.n204 m1m2.n203 0.849769
R5271 m1m2.n205 m1m2.n204 0.849769
R5272 m1m2.n206 m1m2.n205 0.849769
R5273 m1m2.n207 m1m2.n206 0.849769
R5274 m1m2.n208 m1m2.n207 0.849769
R5275 m1m2.n209 m1m2.n208 0.849769
R5276 m1m2.n210 m1m2.n209 0.849769
R5277 m1m2.n211 m1m2.n210 0.849769
R5278 m1m2.n212 m1m2.n211 0.849769
R5279 m1m2.n213 m1m2.n212 0.849769
R5280 m1m2.n214 m1m2.n213 0.849769
R5281 m1m2.n215 m1m2.n214 0.849769
R5282 m1m2.n216 m1m2.n215 0.849769
R5283 m1m2.n217 m1m2.n216 0.849769
R5284 m1m2.n218 m1m2.n217 0.849769
R5285 m1m2.n219 m1m2.n218 0.849769
R5286 m1m2.n220 m1m2.n219 0.849769
R5287 m1m2.n221 m1m2.n220 0.849769
R5288 m1m2.n222 m1m2.n221 0.849769
R5289 m1m2.n223 m1m2.n222 0.849769
R5290 m1m2.n224 m1m2.n223 0.849769
R5291 m1m2.n225 m1m2.n224 0.849769
R5292 m1m2.n226 m1m2.n225 0.849769
R5293 m1m2.n227 m1m2.n226 0.849769
R5294 m1m2.n228 m1m2.n227 0.849769
R5295 m1m2.n229 m1m2.n228 0.849769
R5296 m1m2.n230 m1m2.n229 0.849769
R5297 m1m2.n231 m1m2.n230 0.849769
R5298 m1m2.n232 m1m2.n231 0.849769
R5299 m1m2.n233 m1m2.n232 0.849769
R5300 m1m2.n234 m1m2.n233 0.849769
R5301 m1m2.n235 m1m2.n234 0.849769
R5302 m1m2.n236 m1m2.n235 0.849769
R5303 m1m2.n237 m1m2.n236 0.849769
R5304 m1m2.n238 m1m2.n237 0.849769
R5305 m1m2.n239 m1m2.n238 0.849769
R5306 m1m2.n240 m1m2.n239 0.849769
R5307 m1m2.n241 m1m2.n240 0.849769
R5308 m1m2.n242 m1m2.n241 0.849769
R5309 m1m2.n243 m1m2.n242 0.849769
R5310 m1m2.n244 m1m2.n243 0.849769
R5311 m1m2.n245 m1m2.n244 0.849769
R5312 m1m2.n246 m1m2.n245 0.849769
R5313 m1m2.n247 m1m2.n246 0.849769
R5314 m1m2.n248 m1m2.n247 0.849769
R5315 m1m2.n249 m1m2.n248 0.849769
R5316 m1m2.n250 m1m2.n249 0.849769
R5317 m1m2.n251 m1m2.n250 0.849769
R5318 m1m2.n252 m1m2.n251 0.849769
R5319 m1m2.n253 m1m2.n252 0.849769
R5320 m1m2.n254 m1m2.n253 0.849769
R5321 m1m2.n255 m1m2.n254 0.849769
R5322 m1m2.n256 m1m2.n255 0.849769
R5323 m1m2.n257 m1m2.n256 0.849769
R5324 m1m2.n258 m1m2.n257 0.849769
R5325 m1m2.n259 m1m2.n258 0.849769
R5326 m1m2.n260 m1m2.n259 0.849769
R5327 m1m2.n261 m1m2.n260 0.849769
R5328 m1m2.n262 m1m2.n261 0.849769
R5329 m1m2.n263 m1m2.n262 0.849769
R5330 m1m2.n264 m1m2.n263 0.849769
R5331 m1m2.n265 m1m2.n264 0.849769
R5332 m1m2.n266 m1m2.n265 0.849769
R5333 m1m2.n267 m1m2.n266 0.849769
R5334 m1m2.n268 m1m2.n267 0.849769
R5335 m1m2.n269 m1m2.n268 0.849769
R5336 m1m2.n270 m1m2.n269 0.849769
R5337 m1m2.n271 m1m2.n270 0.849769
R5338 m1m2.n272 m1m2.n271 0.849769
R5339 m1m2.n273 m1m2.n272 0.849769
R5340 m1m2.n274 m1m2.n273 0.849769
R5341 m1m2.n275 m1m2.n274 0.849769
R5342 m1m2.n276 m1m2.n275 0.849769
R5343 m1m2.n277 m1m2.n276 0.849769
R5344 m1m2.n278 m1m2.n277 0.849769
R5345 m1m2.n279 m1m2.n278 0.849769
R5346 m1m2.n280 m1m2.n279 0.849769
R5347 m1m2.n281 m1m2.n280 0.849769
R5348 m1m2.n282 m1m2.n281 0.849769
R5349 m1m2.n283 m1m2.n282 0.849769
R5350 m1m2.n284 m1m2.n283 0.849769
R5351 m1m2.n285 m1m2.n284 0.849769
R5352 m1m2.n286 m1m2.n285 0.849769
R5353 m1m2.n287 m1m2.n286 0.849769
R5354 m1m2.n288 m1m2.n287 0.849769
R5355 m1m2.n289 m1m2.n288 0.849769
R5356 m1m2.n290 m1m2.n289 0.849769
R5357 m1m2.n291 m1m2.n290 0.849769
R5358 m1m2.n292 m1m2.n291 0.849769
R5359 m1m2.n293 m1m2.n292 0.849769
R5360 m1m2.n294 m1m2.n293 0.849769
R5361 m1m2.n295 m1m2.n294 0.849769
R5362 m1m2.n296 m1m2.n295 0.849769
R5363 m1m2.n100 m1m2.n99 0.849769
R5364 m1m2.n101 m1m2.n100 0.849769
R5365 m1m2.n102 m1m2.n101 0.849769
R5366 m1m2.n103 m1m2.n102 0.849769
R5367 m1m2.n104 m1m2.n103 0.849769
R5368 m1m2.n105 m1m2.n104 0.849769
R5369 m1m2.n106 m1m2.n105 0.849769
R5370 m1m2.n107 m1m2.n106 0.849769
R5371 m1m2.n108 m1m2.n107 0.849769
R5372 m1m2.n109 m1m2.n108 0.849769
R5373 m1m2.n110 m1m2.n109 0.849769
R5374 m1m2.n111 m1m2.n110 0.849769
R5375 m1m2.n112 m1m2.n111 0.849769
R5376 m1m2.n113 m1m2.n112 0.849769
R5377 m1m2.n114 m1m2.n113 0.849769
R5378 m1m2.n115 m1m2.n114 0.849769
R5379 m1m2.n116 m1m2.n115 0.849769
R5380 m1m2.n117 m1m2.n116 0.849769
R5381 m1m2.n118 m1m2.n117 0.849769
R5382 m1m2.n119 m1m2.n118 0.849769
R5383 m1m2.n120 m1m2.n119 0.849769
R5384 m1m2.n121 m1m2.n120 0.849769
R5385 m1m2.n122 m1m2.n121 0.849769
R5386 m1m2.n123 m1m2.n122 0.849769
R5387 m1m2.n124 m1m2.n123 0.849769
R5388 m1m2.n125 m1m2.n124 0.849769
R5389 m1m2.n126 m1m2.n125 0.849769
R5390 m1m2.n127 m1m2.n126 0.849769
R5391 m1m2.n128 m1m2.n127 0.849769
R5392 m1m2.n129 m1m2.n128 0.849769
R5393 m1m2.n130 m1m2.n129 0.849769
R5394 m1m2.n131 m1m2.n130 0.849769
R5395 m1m2.n132 m1m2.n131 0.849769
R5396 m1m2.n133 m1m2.n132 0.849769
R5397 m1m2.n134 m1m2.n133 0.849769
R5398 m1m2.n135 m1m2.n134 0.849769
R5399 m1m2.n136 m1m2.n135 0.849769
R5400 m1m2.n137 m1m2.n136 0.849769
R5401 m1m2.n138 m1m2.n137 0.849769
R5402 m1m2.n139 m1m2.n138 0.849769
R5403 m1m2.n140 m1m2.n139 0.849769
R5404 m1m2.n141 m1m2.n140 0.849769
R5405 m1m2.n142 m1m2.n141 0.849769
R5406 m1m2.n143 m1m2.n142 0.849769
R5407 m1m2.n144 m1m2.n143 0.849769
R5408 m1m2.n145 m1m2.n144 0.849769
R5409 m1m2.n146 m1m2.n145 0.849769
R5410 m1m2.n147 m1m2.n146 0.849769
R5411 m1m2.n148 m1m2.n147 0.849769
R5412 m1m2.n149 m1m2.n148 0.849769
R5413 m1m2.n150 m1m2.n149 0.849769
R5414 m1m2.n151 m1m2.n150 0.849769
R5415 m1m2.n152 m1m2.n151 0.849769
R5416 m1m2.n153 m1m2.n152 0.849769
R5417 m1m2.n154 m1m2.n153 0.849769
R5418 m1m2.n155 m1m2.n154 0.849769
R5419 m1m2.n156 m1m2.n155 0.849769
R5420 m1m2.n157 m1m2.n156 0.849769
R5421 m1m2.n158 m1m2.n157 0.849769
R5422 m1m2.n159 m1m2.n158 0.849769
R5423 m1m2.n160 m1m2.n159 0.849769
R5424 m1m2.n161 m1m2.n160 0.849769
R5425 m1m2.n162 m1m2.n161 0.849769
R5426 m1m2.n163 m1m2.n162 0.849769
R5427 m1m2.n164 m1m2.n163 0.849769
R5428 m1m2.n165 m1m2.n164 0.849769
R5429 m1m2.n166 m1m2.n165 0.849769
R5430 m1m2.n167 m1m2.n166 0.849769
R5431 m1m2.n168 m1m2.n167 0.849769
R5432 m1m2.n169 m1m2.n168 0.849769
R5433 m1m2.n170 m1m2.n169 0.849769
R5434 m1m2.n171 m1m2.n170 0.849769
R5435 m1m2.n172 m1m2.n171 0.849769
R5436 m1m2.n173 m1m2.n172 0.849769
R5437 m1m2.n174 m1m2.n173 0.849769
R5438 m1m2.n175 m1m2.n174 0.849769
R5439 m1m2.n176 m1m2.n175 0.849769
R5440 m1m2.n177 m1m2.n176 0.849769
R5441 m1m2.n178 m1m2.n177 0.849769
R5442 m1m2.n179 m1m2.n178 0.849769
R5443 m1m2.n180 m1m2.n179 0.849769
R5444 m1m2.n181 m1m2.n180 0.849769
R5445 m1m2.n182 m1m2.n181 0.849769
R5446 m1m2.n183 m1m2.n182 0.849769
R5447 m1m2.n184 m1m2.n183 0.849769
R5448 m1m2.n185 m1m2.n184 0.849769
R5449 m1m2.n186 m1m2.n185 0.849769
R5450 m1m2.n187 m1m2.n186 0.849769
R5451 m1m2.n188 m1m2.n187 0.849769
R5452 m1m2.n189 m1m2.n188 0.849769
R5453 m1m2.n190 m1m2.n189 0.849769
R5454 m1m2.n191 m1m2.n190 0.849769
R5455 m1m2.n192 m1m2.n191 0.849769
R5456 m1m2.n193 m1m2.n192 0.849769
R5457 m1m2.n194 m1m2.n193 0.849769
R5458 m1m2.n195 m1m2.n194 0.849769
R5459 m1m2.n196 m1m2.n195 0.849769
R5460 m1m2.n197 m1m2.n196 0.849769
R5461 m1m2.n1 m1m2.n0 0.849769
R5462 m1m2.n2 m1m2.n1 0.849769
R5463 m1m2.n3 m1m2.n2 0.849769
R5464 m1m2.n4 m1m2.n3 0.849769
R5465 m1m2.n5 m1m2.n4 0.849769
R5466 m1m2.n6 m1m2.n5 0.849769
R5467 m1m2.n7 m1m2.n6 0.849769
R5468 m1m2.n8 m1m2.n7 0.849769
R5469 m1m2.n9 m1m2.n8 0.849769
R5470 m1m2.n10 m1m2.n9 0.849769
R5471 m1m2.n11 m1m2.n10 0.849769
R5472 m1m2.n12 m1m2.n11 0.849769
R5473 m1m2.n13 m1m2.n12 0.849769
R5474 m1m2.n14 m1m2.n13 0.849769
R5475 m1m2.n15 m1m2.n14 0.849769
R5476 m1m2.n16 m1m2.n15 0.849769
R5477 m1m2.n17 m1m2.n16 0.849769
R5478 m1m2.n18 m1m2.n17 0.849769
R5479 m1m2.n19 m1m2.n18 0.849769
R5480 m1m2.n20 m1m2.n19 0.849769
R5481 m1m2.n21 m1m2.n20 0.849769
R5482 m1m2.n22 m1m2.n21 0.849769
R5483 m1m2.n23 m1m2.n22 0.849769
R5484 m1m2.n24 m1m2.n23 0.849769
R5485 m1m2.n25 m1m2.n24 0.849769
R5486 m1m2.n26 m1m2.n25 0.849769
R5487 m1m2.n27 m1m2.n26 0.849769
R5488 m1m2.n28 m1m2.n27 0.849769
R5489 m1m2.n29 m1m2.n28 0.849769
R5490 m1m2.n30 m1m2.n29 0.849769
R5491 m1m2.n31 m1m2.n30 0.849769
R5492 m1m2.n32 m1m2.n31 0.849769
R5493 m1m2.n33 m1m2.n32 0.849769
R5494 m1m2.n34 m1m2.n33 0.849769
R5495 m1m2.n35 m1m2.n34 0.849769
R5496 m1m2.n36 m1m2.n35 0.849769
R5497 m1m2.n37 m1m2.n36 0.849769
R5498 m1m2.n38 m1m2.n37 0.849769
R5499 m1m2.n39 m1m2.n38 0.849769
R5500 m1m2.n40 m1m2.n39 0.849769
R5501 m1m2.n41 m1m2.n40 0.849769
R5502 m1m2.n42 m1m2.n41 0.849769
R5503 m1m2.n43 m1m2.n42 0.849769
R5504 m1m2.n44 m1m2.n43 0.849769
R5505 m1m2.n45 m1m2.n44 0.849769
R5506 m1m2.n46 m1m2.n45 0.849769
R5507 m1m2.n47 m1m2.n46 0.849769
R5508 m1m2.n48 m1m2.n47 0.849769
R5509 m1m2.n49 m1m2.n48 0.849769
R5510 m1m2.n50 m1m2.n49 0.849769
R5511 m1m2.n51 m1m2.n50 0.849769
R5512 m1m2.n52 m1m2.n51 0.849769
R5513 m1m2.n53 m1m2.n52 0.849769
R5514 m1m2.n54 m1m2.n53 0.849769
R5515 m1m2.n55 m1m2.n54 0.849769
R5516 m1m2.n56 m1m2.n55 0.849769
R5517 m1m2.n57 m1m2.n56 0.849769
R5518 m1m2.n58 m1m2.n57 0.849769
R5519 m1m2.n59 m1m2.n58 0.849769
R5520 m1m2.n60 m1m2.n59 0.849769
R5521 m1m2.n61 m1m2.n60 0.849769
R5522 m1m2.n62 m1m2.n61 0.849769
R5523 m1m2.n63 m1m2.n62 0.849769
R5524 m1m2.n64 m1m2.n63 0.849769
R5525 m1m2.n65 m1m2.n64 0.849769
R5526 m1m2.n66 m1m2.n65 0.849769
R5527 m1m2.n67 m1m2.n66 0.849769
R5528 m1m2.n68 m1m2.n67 0.849769
R5529 m1m2.n69 m1m2.n68 0.849769
R5530 m1m2.n70 m1m2.n69 0.849769
R5531 m1m2.n71 m1m2.n70 0.849769
R5532 m1m2.n72 m1m2.n71 0.849769
R5533 m1m2.n73 m1m2.n72 0.849769
R5534 m1m2.n74 m1m2.n73 0.849769
R5535 m1m2.n75 m1m2.n74 0.849769
R5536 m1m2.n76 m1m2.n75 0.849769
R5537 m1m2.n77 m1m2.n76 0.849769
R5538 m1m2.n78 m1m2.n77 0.849769
R5539 m1m2.n79 m1m2.n78 0.849769
R5540 m1m2.n494 m1m2.n493 0.849769
R5541 m1m2.n493 m1m2.n492 0.849769
R5542 m1m2.n492 m1m2.n491 0.849769
R5543 m1m2.n491 m1m2.n490 0.849769
R5544 m1m2.n490 m1m2.n489 0.849769
R5545 m1m2.n489 m1m2.n488 0.849769
R5546 m1m2.n488 m1m2.n487 0.849769
R5547 m1m2.n487 m1m2.n486 0.849769
R5548 m1m2.n486 m1m2.n485 0.849769
R5549 m1m2.n485 m1m2.n484 0.849769
R5550 m1m2.n484 m1m2.n483 0.849769
R5551 m1m2.n85 m1m2.n84 0.791187
R5552 m1m2.n91 m1m2.n90 0.791187
R5553 m1m2.n93 m1m2.n92 0.791187
R5554 m1m2.n97 m1m2.n96 0.791187
R5555 m1m2.n84 m1m2.n83 0.786223
R5556 m1m2.n80 m1m2.n79 0.772322
R5557 m1m2.n83 m1m2.n82 0.746506
R5558 m1m2.n81 m1m2.n80 0.741542
R5559 m1m2.n82 m1m2.n81 0.741542
R5560 m1m2.n86 m1m2.n85 0.741542
R5561 m1m2.n88 m1m2.n87 0.741542
R5562 m1m2.n89 m1m2.n88 0.741542
R5563 m1m2.n94 m1m2.n93 0.741542
R5564 m1m2.n95 m1m2.n94 0.741542
R5565 m1m2.n96 m1m2.n95 0.741542
R5566 m1m2.n98 m1m2.n97 0.741542
R5567 m1m2.n87 m1m2.n86 0.741542
R5568 m1m2.n90 m1m2.n89 0.741542
R5569 m1m2.n92 m1m2.n91 0.691896
R5570 m1m2.n500 m1m2.n499 0.40943
R5571 m1m2.n501 m1m2.n500 0.40943
R5572 m1m2.n502 m1m2.n501 0.40943
R5573 m1m2.n503 m1m2.n502 0.40943
R5574 m1m2.n504 m1m2.n503 0.40943
R5575 m1m2.n505 m1m2.n504 0.40943
R5576 m1m2.n506 m1m2.n505 0.40943
R5577 m1m2.n507 m1m2.n506 0.40943
R5578 m1m2.n508 m1m2.n507 0.40943
R5579 m1m2.n509 m1m2.n508 0.40943
R5580 m1m2.n510 m1m2.n509 0.40943
R5581 m1m2.n511 m1m2.n510 0.40943
R5582 m1m2.n512 m1m2.n511 0.40943
R5583 m1m2.n513 m1m2.n512 0.40943
R5584 VB_B.n67 VB_B.t62 13.5734
R5585 VB_B.n50 VB_B.t19 13.5734
R5586 VB_B.n33 VB_B.t84 13.5734
R5587 VB_B.n16 VB_B.t29 13.5734
R5588 VB_B.n84 VB_B.t7 13.573
R5589 VB_B.n0 VB_B.t39 13.573
R5590 VB_B.n84 VB_B.t94 13.3193
R5591 VB_B.n85 VB_B.t99 13.3193
R5592 VB_B.n86 VB_B.t2 13.3193
R5593 VB_B.n87 VB_B.t4 13.3193
R5594 VB_B.n88 VB_B.t90 13.3193
R5595 VB_B.n89 VB_B.t97 13.3193
R5596 VB_B.n90 VB_B.t44 13.3193
R5597 VB_B.n91 VB_B.t49 13.3193
R5598 VB_B.n92 VB_B.t55 13.3193
R5599 VB_B.n93 VB_B.t27 13.3193
R5600 VB_B.n94 VB_B.t38 13.3193
R5601 VB_B.n95 VB_B.t14 13.3193
R5602 VB_B.n96 VB_B.t21 13.3193
R5603 VB_B.n97 VB_B.t32 13.3193
R5604 VB_B.n98 VB_B.t65 13.3193
R5605 VB_B.n99 VB_B.t71 13.3193
R5606 VB_B.n67 VB_B.t6 13.3193
R5607 VB_B.n68 VB_B.t10 13.3193
R5608 VB_B.n69 VB_B.t17 13.3193
R5609 VB_B.n70 VB_B.t24 13.3193
R5610 VB_B.n71 VB_B.t37 13.3193
R5611 VB_B.n72 VB_B.t8 13.3193
R5612 VB_B.n73 VB_B.t63 13.3193
R5613 VB_B.n74 VB_B.t67 13.3193
R5614 VB_B.n75 VB_B.t78 13.3193
R5615 VB_B.n76 VB_B.t85 13.3193
R5616 VB_B.n77 VB_B.t59 13.3193
R5617 VB_B.n78 VB_B.t45 13.3193
R5618 VB_B.n79 VB_B.t50 13.3193
R5619 VB_B.n80 VB_B.t56 13.3193
R5620 VB_B.n81 VB_B.t11 13.3193
R5621 VB_B.n82 VB_B.t93 13.3193
R5622 VB_B.n50 VB_B.t74 13.3193
R5623 VB_B.n51 VB_B.t77 13.3193
R5624 VB_B.n52 VB_B.t82 13.3193
R5625 VB_B.n53 VB_B.t88 13.3193
R5626 VB_B.n54 VB_B.t100 13.3193
R5627 VB_B.n55 VB_B.t76 13.3193
R5628 VB_B.n56 VB_B.t75 13.3193
R5629 VB_B.n57 VB_B.t79 13.3193
R5630 VB_B.n58 VB_B.t91 13.3193
R5631 VB_B.n59 VB_B.t98 13.3193
R5632 VB_B.n60 VB_B.t72 13.3193
R5633 VB_B.n61 VB_B.t53 13.3193
R5634 VB_B.n62 VB_B.t57 13.3193
R5635 VB_B.n63 VB_B.t68 13.3193
R5636 VB_B.n64 VB_B.t25 13.3193
R5637 VB_B.n65 VB_B.t1 13.3193
R5638 VB_B.n33 VB_B.t28 13.3193
R5639 VB_B.n34 VB_B.t40 13.3193
R5640 VB_B.n35 VB_B.t47 13.3193
R5641 VB_B.n36 VB_B.t52 13.3193
R5642 VB_B.n37 VB_B.t60 13.3193
R5643 VB_B.n38 VB_B.t33 13.3193
R5644 VB_B.n39 VB_B.t86 13.3193
R5645 VB_B.n40 VB_B.t92 13.3193
R5646 VB_B.n41 VB_B.t0 13.3193
R5647 VB_B.n42 VB_B.t3 13.3193
R5648 VB_B.n43 VB_B.t81 13.3193
R5649 VB_B.n44 VB_B.t64 13.3193
R5650 VB_B.n45 VB_B.t70 13.3193
R5651 VB_B.n46 VB_B.t80 13.3193
R5652 VB_B.n47 VB_B.t41 13.3193
R5653 VB_B.n48 VB_B.t9 13.3193
R5654 VB_B.n16 VB_B.t83 13.3193
R5655 VB_B.n17 VB_B.t89 13.3193
R5656 VB_B.n18 VB_B.t96 13.3193
R5657 VB_B.n19 VB_B.t101 13.3193
R5658 VB_B.n20 VB_B.t5 13.3193
R5659 VB_B.n21 VB_B.t87 13.3193
R5660 VB_B.n22 VB_B.t42 13.3193
R5661 VB_B.n23 VB_B.t48 13.3193
R5662 VB_B.n24 VB_B.t54 13.3193
R5663 VB_B.n25 VB_B.t61 13.3193
R5664 VB_B.n26 VB_B.t35 13.3193
R5665 VB_B.n27 VB_B.t13 13.3193
R5666 VB_B.n28 VB_B.t20 13.3193
R5667 VB_B.n29 VB_B.t30 13.3193
R5668 VB_B.n30 VB_B.t95 13.3193
R5669 VB_B.n31 VB_B.t69 13.3193
R5670 VB_B.n0 VB_B.t15 13.3193
R5671 VB_B.n1 VB_B.t22 13.3193
R5672 VB_B.n2 VB_B.t26 13.3193
R5673 VB_B.n3 VB_B.t34 13.3193
R5674 VB_B.n4 VB_B.t12 13.3193
R5675 VB_B.n5 VB_B.t18 13.3193
R5676 VB_B.n6 VB_B.t46 13.3193
R5677 VB_B.n7 VB_B.t51 13.3193
R5678 VB_B.n8 VB_B.t58 13.3193
R5679 VB_B.n9 VB_B.t31 13.3193
R5680 VB_B.n10 VB_B.t43 13.3193
R5681 VB_B.n11 VB_B.t16 13.3193
R5682 VB_B.n12 VB_B.t23 13.3193
R5683 VB_B.n13 VB_B.t36 13.3193
R5684 VB_B.n14 VB_B.t66 13.3193
R5685 VB_B.n15 VB_B.t73 13.3193
R5686 VB_B VB_B.n100 2.22546
R5687 VB_B.n32 VB_B.n15 0.639878
R5688 VB_B.n100 VB_B.n83 0.460321
R5689 VB_B.n49 VB_B.n32 0.429071
R5690 VB_B.n66 VB_B.n49 0.429071
R5691 VB_B.n83 VB_B.n66 0.429071
R5692 VB_B.n85 VB_B.n84 0.254255
R5693 VB_B.n86 VB_B.n85 0.254255
R5694 VB_B.n87 VB_B.n86 0.254255
R5695 VB_B.n88 VB_B.n87 0.254255
R5696 VB_B.n89 VB_B.n88 0.254255
R5697 VB_B.n90 VB_B.n89 0.254255
R5698 VB_B.n91 VB_B.n90 0.254255
R5699 VB_B.n92 VB_B.n91 0.254255
R5700 VB_B.n93 VB_B.n92 0.254255
R5701 VB_B.n94 VB_B.n93 0.254255
R5702 VB_B.n95 VB_B.n94 0.254255
R5703 VB_B.n96 VB_B.n95 0.254255
R5704 VB_B.n97 VB_B.n96 0.254255
R5705 VB_B.n98 VB_B.n97 0.254255
R5706 VB_B.n99 VB_B.n98 0.254255
R5707 VB_B.n68 VB_B.n67 0.254255
R5708 VB_B.n69 VB_B.n68 0.254255
R5709 VB_B.n70 VB_B.n69 0.254255
R5710 VB_B.n71 VB_B.n70 0.254255
R5711 VB_B.n72 VB_B.n71 0.254255
R5712 VB_B.n73 VB_B.n72 0.254255
R5713 VB_B.n74 VB_B.n73 0.254255
R5714 VB_B.n75 VB_B.n74 0.254255
R5715 VB_B.n76 VB_B.n75 0.254255
R5716 VB_B.n77 VB_B.n76 0.254255
R5717 VB_B.n78 VB_B.n77 0.254255
R5718 VB_B.n79 VB_B.n78 0.254255
R5719 VB_B.n80 VB_B.n79 0.254255
R5720 VB_B.n81 VB_B.n80 0.254255
R5721 VB_B.n82 VB_B.n81 0.254255
R5722 VB_B.n51 VB_B.n50 0.254255
R5723 VB_B.n52 VB_B.n51 0.254255
R5724 VB_B.n53 VB_B.n52 0.254255
R5725 VB_B.n54 VB_B.n53 0.254255
R5726 VB_B.n55 VB_B.n54 0.254255
R5727 VB_B.n56 VB_B.n55 0.254255
R5728 VB_B.n57 VB_B.n56 0.254255
R5729 VB_B.n58 VB_B.n57 0.254255
R5730 VB_B.n59 VB_B.n58 0.254255
R5731 VB_B.n60 VB_B.n59 0.254255
R5732 VB_B.n61 VB_B.n60 0.254255
R5733 VB_B.n62 VB_B.n61 0.254255
R5734 VB_B.n63 VB_B.n62 0.254255
R5735 VB_B.n64 VB_B.n63 0.254255
R5736 VB_B.n65 VB_B.n64 0.254255
R5737 VB_B.n34 VB_B.n33 0.254255
R5738 VB_B.n35 VB_B.n34 0.254255
R5739 VB_B.n36 VB_B.n35 0.254255
R5740 VB_B.n37 VB_B.n36 0.254255
R5741 VB_B.n38 VB_B.n37 0.254255
R5742 VB_B.n39 VB_B.n38 0.254255
R5743 VB_B.n40 VB_B.n39 0.254255
R5744 VB_B.n41 VB_B.n40 0.254255
R5745 VB_B.n42 VB_B.n41 0.254255
R5746 VB_B.n43 VB_B.n42 0.254255
R5747 VB_B.n44 VB_B.n43 0.254255
R5748 VB_B.n45 VB_B.n44 0.254255
R5749 VB_B.n46 VB_B.n45 0.254255
R5750 VB_B.n47 VB_B.n46 0.254255
R5751 VB_B.n48 VB_B.n47 0.254255
R5752 VB_B.n17 VB_B.n16 0.254255
R5753 VB_B.n18 VB_B.n17 0.254255
R5754 VB_B.n19 VB_B.n18 0.254255
R5755 VB_B.n20 VB_B.n19 0.254255
R5756 VB_B.n21 VB_B.n20 0.254255
R5757 VB_B.n22 VB_B.n21 0.254255
R5758 VB_B.n23 VB_B.n22 0.254255
R5759 VB_B.n24 VB_B.n23 0.254255
R5760 VB_B.n25 VB_B.n24 0.254255
R5761 VB_B.n26 VB_B.n25 0.254255
R5762 VB_B.n27 VB_B.n26 0.254255
R5763 VB_B.n28 VB_B.n27 0.254255
R5764 VB_B.n29 VB_B.n28 0.254255
R5765 VB_B.n30 VB_B.n29 0.254255
R5766 VB_B.n31 VB_B.n30 0.254255
R5767 VB_B.n1 VB_B.n0 0.254255
R5768 VB_B.n2 VB_B.n1 0.254255
R5769 VB_B.n3 VB_B.n2 0.254255
R5770 VB_B.n4 VB_B.n3 0.254255
R5771 VB_B.n5 VB_B.n4 0.254255
R5772 VB_B.n6 VB_B.n5 0.254255
R5773 VB_B.n7 VB_B.n6 0.254255
R5774 VB_B.n8 VB_B.n7 0.254255
R5775 VB_B.n9 VB_B.n8 0.254255
R5776 VB_B.n10 VB_B.n9 0.254255
R5777 VB_B.n11 VB_B.n10 0.254255
R5778 VB_B.n12 VB_B.n11 0.254255
R5779 VB_B.n13 VB_B.n12 0.254255
R5780 VB_B.n14 VB_B.n13 0.254255
R5781 VB_B.n15 VB_B.n14 0.254255
R5782 VB_B.n100 VB_B.n99 0.213836
R5783 VB_B.n83 VB_B.n82 0.213419
R5784 VB_B.n66 VB_B.n65 0.213419
R5785 VB_B.n49 VB_B.n48 0.213419
R5786 VB_B.n32 VB_B.n31 0.213419
R5787 m3m4 m3m4.t30 13.474
R5788 m3m4.n28 m3m4.n27 7.12078
R5789 m3m4.n28 m3m4.n13 5.28748
R5790 m3m4.n14 m3m4.t13 4.44742
R5791 m3m4.n0 m3m4.t26 4.42883
R5792 m3m4.n7 m3m4.t29 3.48118
R5793 m3m4.n8 m3m4.t28 3.48118
R5794 m3m4.n9 m3m4.t7 3.48118
R5795 m3m4.n10 m3m4.t17 3.48118
R5796 m3m4.n11 m3m4.t15 3.48118
R5797 m3m4.n12 m3m4.t8 3.48118
R5798 m3m4.n13 m3m4.t23 3.48118
R5799 m3m4.n27 m3m4.t27 3.48118
R5800 m3m4.n26 m3m4.t16 3.48118
R5801 m3m4.n25 m3m4.t19 3.48118
R5802 m3m4.n24 m3m4.t20 3.48118
R5803 m3m4.n23 m3m4.t14 3.48118
R5804 m3m4.n22 m3m4.t1 3.48118
R5805 m3m4.n21 m3m4.t3 3.48118
R5806 m3m4.n20 m3m4.t9 3.48118
R5807 m3m4.n19 m3m4.t12 3.48118
R5808 m3m4.n18 m3m4.t11 3.48118
R5809 m3m4.n17 m3m4.t0 3.48118
R5810 m3m4.n16 m3m4.t4 3.48118
R5811 m3m4.n15 m3m4.t6 3.48118
R5812 m3m4.n14 m3m4.t10 3.48118
R5813 m3m4.n6 m3m4.t2 3.48118
R5814 m3m4.n5 m3m4.t5 3.48118
R5815 m3m4.n4 m3m4.t25 3.48118
R5816 m3m4.n3 m3m4.t18 3.48118
R5817 m3m4.n2 m3m4.t21 3.48118
R5818 m3m4.n1 m3m4.t22 3.48118
R5819 m3m4.n0 m3m4.t24 3.48118
R5820 m3m4 m3m4.n28 1.94529
R5821 m3m4.n15 m3m4.n14 0.966748
R5822 m3m4.n16 m3m4.n15 0.966748
R5823 m3m4.n17 m3m4.n16 0.966748
R5824 m3m4.n18 m3m4.n17 0.966748
R5825 m3m4.n19 m3m4.n18 0.966748
R5826 m3m4.n20 m3m4.n19 0.966748
R5827 m3m4.n21 m3m4.n20 0.966748
R5828 m3m4.n22 m3m4.n21 0.966748
R5829 m3m4.n23 m3m4.n22 0.966748
R5830 m3m4.n24 m3m4.n23 0.966748
R5831 m3m4.n25 m3m4.n24 0.966748
R5832 m3m4.n26 m3m4.n25 0.966748
R5833 m3m4.n27 m3m4.n26 0.966748
R5834 m3m4.n13 m3m4.n12 0.948155
R5835 m3m4.n12 m3m4.n11 0.948155
R5836 m3m4.n11 m3m4.n10 0.948155
R5837 m3m4.n10 m3m4.n9 0.948155
R5838 m3m4.n9 m3m4.n8 0.948155
R5839 m3m4.n8 m3m4.n7 0.948155
R5840 m3m4.n1 m3m4.n0 0.948155
R5841 m3m4.n2 m3m4.n1 0.948155
R5842 m3m4.n3 m3m4.n2 0.948155
R5843 m3m4.n4 m3m4.n3 0.948155
R5844 m3m4.n5 m3m4.n4 0.948155
R5845 m3m4.n6 m3m4.n5 0.948155
R5846 m3m4.n7 m3m4.n6 0.948155
R5847 VSS.n1 VSS.t6 424.322
R5848 VSS.n8 VSS.n0 246.25
R5849 VSS.n6 VSS.n1 136.448
R5850 VSS.t5 VSS.t7 111.96
R5851 VSS.n4 VSS.t9 91.3273
R5852 VSS.n2 VSS.t5 56.1401
R5853 VSS.t8 VSS.n2 55.8202
R5854 VSS.t9 VSS.t10 39.986
R5855 VSS.t11 VSS.t8 31.9889
R5856 VSS.t10 VSS.t0 30.3894
R5857 VSS.t0 VSS.t2 30.3894
R5858 VSS.t14 VSS.t12 30.3894
R5859 VSS.t12 VSS.t11 30.3894
R5860 VSS.t4 VSS.t14 19.1935
R5861 VSS.n7 VSS.n6 14.7205
R5862 VSS.n8 VSS.n7 14.0805
R5863 VSS.n26 VSS.t18 13.9238
R5864 VSS.n26 VSS.t3 13.9238
R5865 VSS.n29 VSS.t19 13.9238
R5866 VSS.n29 VSS.t16 13.9238
R5867 VSS.n28 VSS.t20 13.9238
R5868 VSS.n28 VSS.t15 13.9238
R5869 VSS.n27 VSS.t21 13.9238
R5870 VSS.n27 VSS.t17 13.9238
R5871 VSS.t2 VSS.t4 11.1964
R5872 VSS.n11 VSS.n9 7.99759
R5873 VSS.n31 VSS.t13 6.59787
R5874 VSS.n32 VSS.t1 5.73077
R5875 VSS.n24 VSS.n23 5.32411
R5876 VSS.n13 VSS.n11 5.32186
R5877 VSS.n33 VSS.n32 5.2505
R5878 VSS.n32 VSS.n31 0.882444
R5879 VSS.n28 VSS.n27 0.436512
R5880 VSS.n29 VSS.n28 0.436512
R5881 VSS.n30 VSS.n29 0.22646
R5882 VSS.n30 VSS.n26 0.210551
R5883 VSS VSS.n34 0.165
R5884 VSS.n34 VSS.n33 0.13445
R5885 VSS.n25 VSS.n24 0.00100016
R5886 VSS.n24 VSS.n20 0.00100016
R5887 VSS.n14 VSS.n13 0.00100001
R5888 VSS.n18 VSS.n17 0.00100001
R5889 VSS.n13 VSS.n12 0.001
R5890 VSS.n17 VSS.n16 0.001
R5891 VSS.n31 VSS.n30 0.000511622
R5892 VSS.n23 VSS.n22 0.000504812
R5893 VSS.n11 VSS.n10 0.000504812
R5894 VSS.n23 VSS.n21 0.000504812
R5895 VSS.n6 VSS.n5 0.000501315
R5896 VSS.n5 VSS.n4 0.000501315
R5897 VSS.n9 VSS.n8 0.00050085
R5898 VSS.n4 VSS.n3 0.000500218
R5899 VSS.n34 VSS.n25 0.000500009
R5900 VSS.n16 VSS.n15 0.000500009
R5901 VSS.n20 VSS.n19 0.000500008
R5902 VSS.n19 VSS.n14 0.000500008
R5903 VSS.n19 VSS.n18 0.000500008
R5904 dummy_9.n348 dummy_9.t275 6.56346
R5905 dummy_9.n6 dummy_9.t420 6.41225
R5906 dummy_9.n346 dummy_9.t441 5.77265
R5907 dummy_9.n344 dummy_9.t103 5.77265
R5908 dummy_9.n342 dummy_9.t221 5.77265
R5909 dummy_9.n340 dummy_9.t141 5.77265
R5910 dummy_9.n338 dummy_9.t255 5.77265
R5911 dummy_9.n336 dummy_9.t5 5.77265
R5912 dummy_9.n334 dummy_9.t307 5.77265
R5913 dummy_9.n332 dummy_9.t439 5.77265
R5914 dummy_9.n330 dummy_9.t351 5.77265
R5915 dummy_9.n328 dummy_9.t35 5.77265
R5916 dummy_9.n347 dummy_9.t440 5.77129
R5917 dummy_9.n345 dummy_9.t102 5.77129
R5918 dummy_9.n343 dummy_9.t220 5.77129
R5919 dummy_9.n341 dummy_9.t140 5.77129
R5920 dummy_9.n339 dummy_9.t254 5.77129
R5921 dummy_9.n337 dummy_9.t4 5.77129
R5922 dummy_9.n335 dummy_9.t306 5.77129
R5923 dummy_9.n333 dummy_9.t438 5.77129
R5924 dummy_9.n331 dummy_9.t350 5.77129
R5925 dummy_9.n329 dummy_9.t34 5.77129
R5926 dummy_9.n327 dummy_9.t184 5.77129
R5927 dummy_9.n127 dummy_9.t279 5.75294
R5928 dummy_9.n107 dummy_9.t151 5.75075
R5929 dummy_9.n109 dummy_9.t197 5.75075
R5930 dummy_9.n111 dummy_9.t161 5.75075
R5931 dummy_9.n113 dummy_9.t205 5.75075
R5932 dummy_9.n115 dummy_9.t11 5.75075
R5933 dummy_9.n117 dummy_9.t223 5.75075
R5934 dummy_9.n119 dummy_9.t263 5.75075
R5935 dummy_9.n121 dummy_9.t235 5.75075
R5936 dummy_9.n123 dummy_9.t283 5.75075
R5937 dummy_9.n125 dummy_9.t325 5.75075
R5938 dummy_9.n108 dummy_9.t150 5.75014
R5939 dummy_9.n110 dummy_9.t196 5.75014
R5940 dummy_9.n112 dummy_9.t160 5.75014
R5941 dummy_9.n114 dummy_9.t204 5.75014
R5942 dummy_9.n116 dummy_9.t10 5.75014
R5943 dummy_9.n118 dummy_9.t222 5.75014
R5944 dummy_9.n120 dummy_9.t262 5.75014
R5945 dummy_9.n122 dummy_9.t234 5.75014
R5946 dummy_9.n124 dummy_9.t282 5.75014
R5947 dummy_9.n126 dummy_9.t324 5.75014
R5948 dummy_9.n326 dummy_9.t185 5.74966
R5949 dummy_9.n447 dummy_9.t130 5.74893
R5950 dummy_9.n0 dummy_9.t131 5.71641
R5951 dummy_9.n105 dummy_9.t214 5.7154
R5952 dummy_9.n5 dummy_9.t215 5.7154
R5953 dummy_9.n128 dummy_9.t278 5.7154
R5954 dummy_9.n370 dummy_9.t273 5.71419
R5955 dummy_9.n369 dummy_9.t165 5.71419
R5956 dummy_9.n368 dummy_9.t285 5.71419
R5957 dummy_9.n367 dummy_9.t393 5.71419
R5958 dummy_9.n366 dummy_9.t257 5.71419
R5959 dummy_9.n365 dummy_9.t379 5.71419
R5960 dummy_9.n364 dummy_9.t153 5.71419
R5961 dummy_9.n363 dummy_9.t387 5.71419
R5962 dummy_9.n362 dummy_9.t237 5.71419
R5963 dummy_9.n361 dummy_9.t29 5.71419
R5964 dummy_9.n360 dummy_9.t227 5.71419
R5965 dummy_9.n359 dummy_9.t39 5.71419
R5966 dummy_9.n358 dummy_9.t233 5.71419
R5967 dummy_9.n357 dummy_9.t317 5.71419
R5968 dummy_9.n356 dummy_9.t115 5.71419
R5969 dummy_9.n355 dummy_9.t329 5.71419
R5970 dummy_9.n354 dummy_9.t331 5.71419
R5971 dummy_9.n353 dummy_9.t423 5.71419
R5972 dummy_9.n352 dummy_9.t167 5.71419
R5973 dummy_9.n351 dummy_9.t431 5.71419
R5974 dummy_9.n350 dummy_9.t85 5.71419
R5975 dummy_9.n349 dummy_9.t407 5.71419
R5976 dummy_9.n348 dummy_9.t79 5.71419
R5977 dummy_9.n372 dummy_9.t179 5.71419
R5978 dummy_9.n373 dummy_9.t435 5.71419
R5979 dummy_9.n374 dummy_9.t313 5.71419
R5980 dummy_9.n375 dummy_9.t7 5.71419
R5981 dummy_9.n376 dummy_9.t339 5.71419
R5982 dummy_9.n377 dummy_9.t93 5.71419
R5983 dummy_9.n378 dummy_9.t327 5.71419
R5984 dummy_9.n379 dummy_9.t225 5.71419
R5985 dummy_9.n380 dummy_9.t3 5.71419
R5986 dummy_9.n381 dummy_9.t217 5.71419
R5987 dummy_9.n382 dummy_9.t443 5.71419
R5988 dummy_9.n383 dummy_9.t321 5.71419
R5989 dummy_9.n384 dummy_9.t133 5.71419
R5990 dummy_9.n385 dummy_9.t341 5.71419
R5991 dummy_9.n386 dummy_9.t129 5.71419
R5992 dummy_9.n387 dummy_9.t337 5.71419
R5993 dummy_9.n388 dummy_9.t55 5.71419
R5994 dummy_9.n389 dummy_9.t271 5.71419
R5995 dummy_9.n390 dummy_9.t45 5.71419
R5996 dummy_9.n391 dummy_9.t383 5.71419
R5997 dummy_9.n392 dummy_9.t63 5.71419
R5998 dummy_9.n393 dummy_9.t397 5.71419
R5999 dummy_9.n394 dummy_9.t287 5.71419
R6000 dummy_9.n395 dummy_9.t391 5.71419
R6001 dummy_9.n396 dummy_9.t91 5.71419
R6002 dummy_9.n397 dummy_9.t299 5.71419
R6003 dummy_9.n398 dummy_9.t87 5.71419
R6004 dummy_9.n399 dummy_9.t437 5.71419
R6005 dummy_9.n400 dummy_9.t97 5.71419
R6006 dummy_9.n401 dummy_9.t15 5.71419
R6007 dummy_9.n402 dummy_9.t191 5.71419
R6008 dummy_9.n403 dummy_9.t1 5.71419
R6009 dummy_9.n404 dummy_9.t125 5.71419
R6010 dummy_9.n405 dummy_9.t355 5.71419
R6011 dummy_9.n406 dummy_9.t137 5.71419
R6012 dummy_9.n407 dummy_9.t347 5.71419
R6013 dummy_9.n408 dummy_9.t231 5.71419
R6014 dummy_9.n409 dummy_9.t59 5.71419
R6015 dummy_9.n410 dummy_9.t239 5.71419
R6016 dummy_9.n411 dummy_9.t53 5.71419
R6017 dummy_9.n412 dummy_9.t51 5.71419
R6018 dummy_9.n413 dummy_9.t405 5.71419
R6019 dummy_9.n414 dummy_9.t175 5.71419
R6020 dummy_9.n415 dummy_9.t399 5.71419
R6021 dummy_9.n416 dummy_9.t291 5.71419
R6022 dummy_9.n417 dummy_9.t419 5.71419
R6023 dummy_9.n418 dummy_9.t305 5.71419
R6024 dummy_9.n419 dummy_9.t187 5.71419
R6025 dummy_9.n420 dummy_9.t89 5.71419
R6026 dummy_9.n421 dummy_9.t445 5.71419
R6027 dummy_9.n422 dummy_9.t203 5.71419
R6028 dummy_9.n423 dummy_9.t17 5.71419
R6029 dummy_9.n424 dummy_9.t343 5.71419
R6030 dummy_9.n425 dummy_9.t9 5.71419
R6031 dummy_9.n426 dummy_9.t363 5.71419
R6032 dummy_9.n427 dummy_9.t119 5.71419
R6033 dummy_9.n428 dummy_9.t139 5.71419
R6034 dummy_9.n429 dummy_9.t47 5.71419
R6035 dummy_9.n430 dummy_9.t249 5.71419
R6036 dummy_9.n431 dummy_9.t67 5.71419
R6037 dummy_9.n432 dummy_9.t243 5.71419
R6038 dummy_9.n433 dummy_9.t145 5.71419
R6039 dummy_9.n434 dummy_9.t413 5.71419
R6040 dummy_9.n435 dummy_9.t155 5.71419
R6041 dummy_9.n436 dummy_9.t183 5.71419
R6042 dummy_9.n437 dummy_9.t403 5.71419
R6043 dummy_9.n438 dummy_9.t295 5.71419
R6044 dummy_9.n439 dummy_9.t101 5.71419
R6045 dummy_9.n440 dummy_9.t309 5.71419
R6046 dummy_9.n441 dummy_9.t193 5.71419
R6047 dummy_9.n442 dummy_9.t301 5.71419
R6048 dummy_9.n443 dummy_9.t209 5.71419
R6049 dummy_9.n444 dummy_9.t359 5.71419
R6050 dummy_9.n445 dummy_9.t21 5.71419
R6051 dummy_9.n446 dummy_9.t349 5.71419
R6052 dummy_9.n228 dummy_9.t348 5.71419
R6053 dummy_9.n227 dummy_9.t20 5.71419
R6054 dummy_9.n226 dummy_9.t358 5.71419
R6055 dummy_9.n225 dummy_9.t208 5.71419
R6056 dummy_9.n224 dummy_9.t300 5.71419
R6057 dummy_9.n223 dummy_9.t192 5.71419
R6058 dummy_9.n222 dummy_9.t308 5.71419
R6059 dummy_9.n221 dummy_9.t100 5.71419
R6060 dummy_9.n220 dummy_9.t294 5.71419
R6061 dummy_9.n219 dummy_9.t402 5.71419
R6062 dummy_9.n218 dummy_9.t182 5.71419
R6063 dummy_9.n217 dummy_9.t154 5.71419
R6064 dummy_9.n216 dummy_9.t412 5.71419
R6065 dummy_9.n215 dummy_9.t144 5.71419
R6066 dummy_9.n214 dummy_9.t242 5.71419
R6067 dummy_9.n213 dummy_9.t66 5.71419
R6068 dummy_9.n212 dummy_9.t248 5.71419
R6069 dummy_9.n211 dummy_9.t46 5.71419
R6070 dummy_9.n210 dummy_9.t138 5.71419
R6071 dummy_9.n209 dummy_9.t118 5.71419
R6072 dummy_9.n208 dummy_9.t362 5.71419
R6073 dummy_9.n207 dummy_9.t8 5.71419
R6074 dummy_9.n206 dummy_9.t342 5.71419
R6075 dummy_9.n205 dummy_9.t16 5.71419
R6076 dummy_9.n204 dummy_9.t202 5.71419
R6077 dummy_9.n203 dummy_9.t444 5.71419
R6078 dummy_9.n202 dummy_9.t88 5.71419
R6079 dummy_9.n201 dummy_9.t186 5.71419
R6080 dummy_9.n200 dummy_9.t304 5.71419
R6081 dummy_9.n199 dummy_9.t418 5.71419
R6082 dummy_9.n198 dummy_9.t290 5.71419
R6083 dummy_9.n197 dummy_9.t398 5.71419
R6084 dummy_9.n196 dummy_9.t174 5.71419
R6085 dummy_9.n195 dummy_9.t404 5.71419
R6086 dummy_9.n194 dummy_9.t50 5.71419
R6087 dummy_9.n193 dummy_9.t52 5.71419
R6088 dummy_9.n192 dummy_9.t238 5.71419
R6089 dummy_9.n191 dummy_9.t58 5.71419
R6090 dummy_9.n190 dummy_9.t230 5.71419
R6091 dummy_9.n189 dummy_9.t346 5.71419
R6092 dummy_9.n188 dummy_9.t136 5.71419
R6093 dummy_9.n187 dummy_9.t354 5.71419
R6094 dummy_9.n186 dummy_9.t124 5.71419
R6095 dummy_9.n185 dummy_9.t0 5.71419
R6096 dummy_9.n184 dummy_9.t190 5.71419
R6097 dummy_9.n183 dummy_9.t14 5.71419
R6098 dummy_9.n182 dummy_9.t96 5.71419
R6099 dummy_9.n181 dummy_9.t436 5.71419
R6100 dummy_9.n180 dummy_9.t86 5.71419
R6101 dummy_9.n179 dummy_9.t298 5.71419
R6102 dummy_9.n178 dummy_9.t90 5.71419
R6103 dummy_9.n177 dummy_9.t390 5.71419
R6104 dummy_9.n176 dummy_9.t286 5.71419
R6105 dummy_9.n175 dummy_9.t396 5.71419
R6106 dummy_9.n174 dummy_9.t62 5.71419
R6107 dummy_9.n173 dummy_9.t382 5.71419
R6108 dummy_9.n172 dummy_9.t44 5.71419
R6109 dummy_9.n171 dummy_9.t270 5.71419
R6110 dummy_9.n170 dummy_9.t54 5.71419
R6111 dummy_9.n169 dummy_9.t336 5.71419
R6112 dummy_9.n168 dummy_9.t128 5.71419
R6113 dummy_9.n167 dummy_9.t340 5.71419
R6114 dummy_9.n166 dummy_9.t132 5.71419
R6115 dummy_9.n165 dummy_9.t320 5.71419
R6116 dummy_9.n164 dummy_9.t442 5.71419
R6117 dummy_9.n163 dummy_9.t216 5.71419
R6118 dummy_9.n162 dummy_9.t2 5.71419
R6119 dummy_9.n161 dummy_9.t224 5.71419
R6120 dummy_9.n160 dummy_9.t326 5.71419
R6121 dummy_9.n159 dummy_9.t92 5.71419
R6122 dummy_9.n158 dummy_9.t338 5.71419
R6123 dummy_9.n157 dummy_9.t6 5.71419
R6124 dummy_9.n156 dummy_9.t312 5.71419
R6125 dummy_9.n155 dummy_9.t434 5.71419
R6126 dummy_9.n154 dummy_9.t178 5.71419
R6127 dummy_9.n153 dummy_9.t446 5.71419
R6128 dummy_9.n152 dummy_9.t272 5.71419
R6129 dummy_9.n151 dummy_9.t164 5.71419
R6130 dummy_9.n150 dummy_9.t284 5.71419
R6131 dummy_9.n149 dummy_9.t392 5.71419
R6132 dummy_9.n148 dummy_9.t256 5.71419
R6133 dummy_9.n147 dummy_9.t378 5.71419
R6134 dummy_9.n146 dummy_9.t152 5.71419
R6135 dummy_9.n145 dummy_9.t386 5.71419
R6136 dummy_9.n144 dummy_9.t236 5.71419
R6137 dummy_9.n143 dummy_9.t28 5.71419
R6138 dummy_9.n142 dummy_9.t226 5.71419
R6139 dummy_9.n141 dummy_9.t38 5.71419
R6140 dummy_9.n140 dummy_9.t232 5.71419
R6141 dummy_9.n139 dummy_9.t316 5.71419
R6142 dummy_9.n138 dummy_9.t114 5.71419
R6143 dummy_9.n137 dummy_9.t328 5.71419
R6144 dummy_9.n136 dummy_9.t330 5.71419
R6145 dummy_9.n135 dummy_9.t422 5.71419
R6146 dummy_9.n134 dummy_9.t166 5.71419
R6147 dummy_9.n133 dummy_9.t430 5.71419
R6148 dummy_9.n132 dummy_9.t84 5.71419
R6149 dummy_9.n131 dummy_9.t406 5.71419
R6150 dummy_9.n130 dummy_9.t78 5.71419
R6151 dummy_9.n129 dummy_9.t274 5.71419
R6152 dummy_9.n104 dummy_9.t212 5.71419
R6153 dummy_9.n103 dummy_9.t22 5.71419
R6154 dummy_9.n102 dummy_9.t352 5.71419
R6155 dummy_9.n101 dummy_9.t36 5.71419
R6156 dummy_9.n100 dummy_9.t368 5.71419
R6157 dummy_9.n99 dummy_9.t126 5.71419
R6158 dummy_9.n98 dummy_9.t364 5.71419
R6159 dummy_9.n97 dummy_9.t268 5.71419
R6160 dummy_9.n96 dummy_9.t266 5.71419
R6161 dummy_9.n95 dummy_9.t72 5.71419
R6162 dummy_9.n94 dummy_9.t252 5.71419
R6163 dummy_9.n93 dummy_9.t168 5.71419
R6164 dummy_9.n92 dummy_9.t424 5.71419
R6165 dummy_9.n91 dummy_9.t162 5.71419
R6166 dummy_9.n90 dummy_9.t414 5.71419
R6167 dummy_9.n89 dummy_9.t176 5.71419
R6168 dummy_9.n88 dummy_9.t318 5.71419
R6169 dummy_9.n87 dummy_9.t110 5.71419
R6170 dummy_9.n86 dummy_9.t310 5.71419
R6171 dummy_9.n85 dummy_9.t200 5.71419
R6172 dummy_9.n84 dummy_9.t334 5.71419
R6173 dummy_9.n83 dummy_9.t218 5.71419
R6174 dummy_9.n82 dummy_9.t122 5.71419
R6175 dummy_9.n81 dummy_9.t210 5.71419
R6176 dummy_9.n80 dummy_9.t380 5.71419
R6177 dummy_9.n79 dummy_9.t134 5.71419
R6178 dummy_9.n78 dummy_9.t372 5.71419
R6179 dummy_9.n77 dummy_9.t246 5.71419
R6180 dummy_9.n76 dummy_9.t388 5.71419
R6181 dummy_9.n75 dummy_9.t276 5.71419
R6182 dummy_9.n74 dummy_9.t48 5.71419
R6183 dummy_9.n73 dummy_9.t264 5.71419
R6184 dummy_9.n72 dummy_9.t296 5.71419
R6185 dummy_9.n71 dummy_9.t70 5.71419
R6186 dummy_9.n70 dummy_9.t292 5.71419
R6187 dummy_9.n69 dummy_9.t60 5.71419
R6188 dummy_9.n68 dummy_9.t394 5.71419
R6189 dummy_9.n67 dummy_9.t188 5.71419
R6190 dummy_9.n66 dummy_9.t408 5.71419
R6191 dummy_9.n65 dummy_9.t180 5.71419
R6192 dummy_9.n64 dummy_9.t400 5.71419
R6193 dummy_9.n63 dummy_9.t108 5.71419
R6194 dummy_9.n62 dummy_9.t344 5.71419
R6195 dummy_9.n61 dummy_9.t94 5.71419
R6196 dummy_9.n60 dummy_9.t12 5.71419
R6197 dummy_9.n59 dummy_9.t116 5.71419
R6198 dummy_9.n58 dummy_9.t24 5.71419
R6199 dummy_9.n57 dummy_9.t356 5.71419
R6200 dummy_9.n56 dummy_9.t18 5.71419
R6201 dummy_9.n55 dummy_9.t148 5.71419
R6202 dummy_9.n54 dummy_9.t370 5.71419
R6203 dummy_9.n53 dummy_9.t142 5.71419
R6204 dummy_9.n52 dummy_9.t56 5.71419
R6205 dummy_9.n51 dummy_9.t156 5.71419
R6206 dummy_9.n50 dummy_9.t76 5.71419
R6207 dummy_9.n49 dummy_9.t258 5.71419
R6208 dummy_9.n48 dummy_9.t68 5.71419
R6209 dummy_9.n47 dummy_9.t172 5.71419
R6210 dummy_9.n46 dummy_9.t426 5.71419
R6211 dummy_9.n45 dummy_9.t194 5.71419
R6212 dummy_9.n44 dummy_9.t416 5.71419
R6213 dummy_9.n43 dummy_9.t302 5.71419
R6214 dummy_9.n42 dummy_9.t112 5.71419
R6215 dummy_9.n41 dummy_9.t314 5.71419
R6216 dummy_9.n40 dummy_9.t106 5.71419
R6217 dummy_9.n39 dummy_9.t104 5.71419
R6218 dummy_9.n38 dummy_9.t32 5.71419
R6219 dummy_9.n37 dummy_9.t240 5.71419
R6220 dummy_9.n36 dummy_9.t26 5.71419
R6221 dummy_9.n35 dummy_9.t360 5.71419
R6222 dummy_9.n34 dummy_9.t42 5.71419
R6223 dummy_9.n33 dummy_9.t376 5.71419
R6224 dummy_9.n32 dummy_9.t250 5.71419
R6225 dummy_9.n31 dummy_9.t146 5.71419
R6226 dummy_9.n30 dummy_9.t64 5.71419
R6227 dummy_9.n29 dummy_9.t280 5.71419
R6228 dummy_9.n28 dummy_9.t80 5.71419
R6229 dummy_9.n27 dummy_9.t410 5.71419
R6230 dummy_9.n26 dummy_9.t74 5.71419
R6231 dummy_9.n25 dummy_9.t432 5.71419
R6232 dummy_9.n24 dummy_9.t170 5.71419
R6233 dummy_9.n23 dummy_9.t198 5.71419
R6234 dummy_9.n22 dummy_9.t98 5.71419
R6235 dummy_9.n21 dummy_9.t332 5.71419
R6236 dummy_9.n20 dummy_9.t120 5.71419
R6237 dummy_9.n19 dummy_9.t322 5.71419
R6238 dummy_9.n18 dummy_9.t206 5.71419
R6239 dummy_9.n17 dummy_9.t40 5.71419
R6240 dummy_9.n16 dummy_9.t228 5.71419
R6241 dummy_9.n15 dummy_9.t244 5.71419
R6242 dummy_9.n14 dummy_9.t30 5.71419
R6243 dummy_9.n13 dummy_9.t366 5.71419
R6244 dummy_9.n12 dummy_9.t158 5.71419
R6245 dummy_9.n11 dummy_9.t384 5.71419
R6246 dummy_9.n10 dummy_9.t260 5.71419
R6247 dummy_9.n9 dummy_9.t374 5.71419
R6248 dummy_9.n8 dummy_9.t288 5.71419
R6249 dummy_9.n7 dummy_9.t428 5.71419
R6250 dummy_9.n6 dummy_9.t82 5.71419
R6251 dummy_9.n4 dummy_9.t213 5.71419
R6252 dummy_9.n3 dummy_9.t23 5.71419
R6253 dummy_9.n2 dummy_9.t353 5.71419
R6254 dummy_9.n229 dummy_9.t37 5.71419
R6255 dummy_9.n230 dummy_9.t369 5.71419
R6256 dummy_9.n231 dummy_9.t127 5.71419
R6257 dummy_9.n232 dummy_9.t365 5.71419
R6258 dummy_9.n233 dummy_9.t269 5.71419
R6259 dummy_9.n234 dummy_9.t267 5.71419
R6260 dummy_9.n235 dummy_9.t73 5.71419
R6261 dummy_9.n236 dummy_9.t253 5.71419
R6262 dummy_9.n237 dummy_9.t169 5.71419
R6263 dummy_9.n238 dummy_9.t425 5.71419
R6264 dummy_9.n239 dummy_9.t163 5.71419
R6265 dummy_9.n240 dummy_9.t415 5.71419
R6266 dummy_9.n241 dummy_9.t177 5.71419
R6267 dummy_9.n242 dummy_9.t319 5.71419
R6268 dummy_9.n243 dummy_9.t111 5.71419
R6269 dummy_9.n244 dummy_9.t311 5.71419
R6270 dummy_9.n245 dummy_9.t201 5.71419
R6271 dummy_9.n246 dummy_9.t335 5.71419
R6272 dummy_9.n247 dummy_9.t219 5.71419
R6273 dummy_9.n248 dummy_9.t123 5.71419
R6274 dummy_9.n249 dummy_9.t211 5.71419
R6275 dummy_9.n250 dummy_9.t381 5.71419
R6276 dummy_9.n251 dummy_9.t135 5.71419
R6277 dummy_9.n252 dummy_9.t373 5.71419
R6278 dummy_9.n253 dummy_9.t247 5.71419
R6279 dummy_9.n254 dummy_9.t389 5.71419
R6280 dummy_9.n255 dummy_9.t277 5.71419
R6281 dummy_9.n256 dummy_9.t49 5.71419
R6282 dummy_9.n257 dummy_9.t265 5.71419
R6283 dummy_9.n258 dummy_9.t297 5.71419
R6284 dummy_9.n259 dummy_9.t71 5.71419
R6285 dummy_9.n260 dummy_9.t293 5.71419
R6286 dummy_9.n261 dummy_9.t61 5.71419
R6287 dummy_9.n262 dummy_9.t395 5.71419
R6288 dummy_9.n263 dummy_9.t189 5.71419
R6289 dummy_9.n264 dummy_9.t409 5.71419
R6290 dummy_9.n265 dummy_9.t181 5.71419
R6291 dummy_9.n266 dummy_9.t401 5.71419
R6292 dummy_9.n267 dummy_9.t109 5.71419
R6293 dummy_9.n268 dummy_9.t345 5.71419
R6294 dummy_9.n269 dummy_9.t95 5.71419
R6295 dummy_9.n270 dummy_9.t13 5.71419
R6296 dummy_9.n271 dummy_9.t117 5.71419
R6297 dummy_9.n272 dummy_9.t25 5.71419
R6298 dummy_9.n273 dummy_9.t357 5.71419
R6299 dummy_9.n274 dummy_9.t19 5.71419
R6300 dummy_9.n275 dummy_9.t149 5.71419
R6301 dummy_9.n276 dummy_9.t371 5.71419
R6302 dummy_9.n277 dummy_9.t143 5.71419
R6303 dummy_9.n278 dummy_9.t57 5.71419
R6304 dummy_9.n279 dummy_9.t157 5.71419
R6305 dummy_9.n280 dummy_9.t77 5.71419
R6306 dummy_9.n281 dummy_9.t259 5.71419
R6307 dummy_9.n282 dummy_9.t69 5.71419
R6308 dummy_9.n283 dummy_9.t173 5.71419
R6309 dummy_9.n284 dummy_9.t427 5.71419
R6310 dummy_9.n285 dummy_9.t195 5.71419
R6311 dummy_9.n286 dummy_9.t417 5.71419
R6312 dummy_9.n287 dummy_9.t303 5.71419
R6313 dummy_9.n288 dummy_9.t113 5.71419
R6314 dummy_9.n289 dummy_9.t315 5.71419
R6315 dummy_9.n290 dummy_9.t107 5.71419
R6316 dummy_9.n291 dummy_9.t105 5.71419
R6317 dummy_9.n292 dummy_9.t33 5.71419
R6318 dummy_9.n293 dummy_9.t241 5.71419
R6319 dummy_9.n294 dummy_9.t27 5.71419
R6320 dummy_9.n295 dummy_9.t361 5.71419
R6321 dummy_9.n296 dummy_9.t43 5.71419
R6322 dummy_9.n297 dummy_9.t377 5.71419
R6323 dummy_9.n298 dummy_9.t251 5.71419
R6324 dummy_9.n299 dummy_9.t147 5.71419
R6325 dummy_9.n300 dummy_9.t65 5.71419
R6326 dummy_9.n301 dummy_9.t281 5.71419
R6327 dummy_9.n302 dummy_9.t81 5.71419
R6328 dummy_9.n303 dummy_9.t411 5.71419
R6329 dummy_9.n304 dummy_9.t75 5.71419
R6330 dummy_9.n305 dummy_9.t433 5.71419
R6331 dummy_9.n306 dummy_9.t171 5.71419
R6332 dummy_9.n307 dummy_9.t199 5.71419
R6333 dummy_9.n308 dummy_9.t99 5.71419
R6334 dummy_9.n309 dummy_9.t333 5.71419
R6335 dummy_9.n310 dummy_9.t121 5.71419
R6336 dummy_9.n311 dummy_9.t323 5.71419
R6337 dummy_9.n312 dummy_9.t207 5.71419
R6338 dummy_9.n313 dummy_9.t41 5.71419
R6339 dummy_9.n314 dummy_9.t229 5.71419
R6340 dummy_9.n315 dummy_9.t245 5.71419
R6341 dummy_9.n316 dummy_9.t31 5.71419
R6342 dummy_9.n317 dummy_9.t367 5.71419
R6343 dummy_9.n318 dummy_9.t159 5.71419
R6344 dummy_9.n319 dummy_9.t385 5.71419
R6345 dummy_9.n320 dummy_9.t261 5.71419
R6346 dummy_9.n321 dummy_9.t375 5.71419
R6347 dummy_9.n322 dummy_9.t289 5.71419
R6348 dummy_9.n323 dummy_9.t429 5.71419
R6349 dummy_9.n324 dummy_9.t83 5.71419
R6350 dummy_9.n325 dummy_9.t421 5.71419
R6351 dummy_9.n371 dummy_9.t447 5.71419
R6352 dummy_9.n447 dummy_9.n0 1.80275
R6353 dummy_9.n106 dummy_9.n5 1.80136
R6354 dummy_9.n128 dummy_9.n127 1.8007
R6355 dummy_9.n327 dummy_9.n326 1.77926
R6356 dummy_9.n347 dummy_9.n346 1.77826
R6357 dummy_9.n345 dummy_9.n344 1.77826
R6358 dummy_9.n343 dummy_9.n342 1.77826
R6359 dummy_9.n341 dummy_9.n340 1.77826
R6360 dummy_9.n339 dummy_9.n338 1.77826
R6361 dummy_9.n337 dummy_9.n336 1.77826
R6362 dummy_9.n335 dummy_9.n334 1.77826
R6363 dummy_9.n333 dummy_9.n332 1.77826
R6364 dummy_9.n331 dummy_9.n330 1.77826
R6365 dummy_9.n329 dummy_9.n328 1.77826
R6366 dummy_9.n126 dummy_9.n125 1.77826
R6367 dummy_9.n124 dummy_9.n123 1.77826
R6368 dummy_9.n122 dummy_9.n121 1.77826
R6369 dummy_9.n120 dummy_9.n119 1.77826
R6370 dummy_9.n118 dummy_9.n117 1.77826
R6371 dummy_9.n116 dummy_9.n115 1.77826
R6372 dummy_9.n114 dummy_9.n113 1.77826
R6373 dummy_9.n112 dummy_9.n111 1.77826
R6374 dummy_9.n110 dummy_9.n109 1.77826
R6375 dummy_9.n108 dummy_9.n107 1.77826
R6376 dummy_9.n1 dummy_9.n446 1.22605
R6377 dummy_9.n349 dummy_9.n348 0.849769
R6378 dummy_9.n350 dummy_9.n349 0.849769
R6379 dummy_9.n351 dummy_9.n350 0.849769
R6380 dummy_9.n352 dummy_9.n351 0.849769
R6381 dummy_9.n353 dummy_9.n352 0.849769
R6382 dummy_9.n354 dummy_9.n353 0.849769
R6383 dummy_9.n355 dummy_9.n354 0.849769
R6384 dummy_9.n356 dummy_9.n355 0.849769
R6385 dummy_9.n357 dummy_9.n356 0.849769
R6386 dummy_9.n358 dummy_9.n357 0.849769
R6387 dummy_9.n359 dummy_9.n358 0.849769
R6388 dummy_9.n360 dummy_9.n359 0.849769
R6389 dummy_9.n361 dummy_9.n360 0.849769
R6390 dummy_9.n362 dummy_9.n361 0.849769
R6391 dummy_9.n363 dummy_9.n362 0.849769
R6392 dummy_9.n364 dummy_9.n363 0.849769
R6393 dummy_9.n365 dummy_9.n364 0.849769
R6394 dummy_9.n366 dummy_9.n365 0.849769
R6395 dummy_9.n367 dummy_9.n366 0.849769
R6396 dummy_9.n368 dummy_9.n367 0.849769
R6397 dummy_9.n369 dummy_9.n368 0.849769
R6398 dummy_9.n370 dummy_9.n369 0.849769
R6399 dummy_9.n371 dummy_9.n370 0.849769
R6400 dummy_9.n325 dummy_9.n324 0.849769
R6401 dummy_9.n324 dummy_9.n323 0.849769
R6402 dummy_9.n323 dummy_9.n322 0.849769
R6403 dummy_9.n322 dummy_9.n321 0.849769
R6404 dummy_9.n321 dummy_9.n320 0.849769
R6405 dummy_9.n320 dummy_9.n319 0.849769
R6406 dummy_9.n319 dummy_9.n318 0.849769
R6407 dummy_9.n318 dummy_9.n317 0.849769
R6408 dummy_9.n317 dummy_9.n316 0.849769
R6409 dummy_9.n316 dummy_9.n315 0.849769
R6410 dummy_9.n315 dummy_9.n314 0.849769
R6411 dummy_9.n314 dummy_9.n313 0.849769
R6412 dummy_9.n313 dummy_9.n312 0.849769
R6413 dummy_9.n312 dummy_9.n311 0.849769
R6414 dummy_9.n311 dummy_9.n310 0.849769
R6415 dummy_9.n310 dummy_9.n309 0.849769
R6416 dummy_9.n309 dummy_9.n308 0.849769
R6417 dummy_9.n308 dummy_9.n307 0.849769
R6418 dummy_9.n307 dummy_9.n306 0.849769
R6419 dummy_9.n306 dummy_9.n305 0.849769
R6420 dummy_9.n305 dummy_9.n304 0.849769
R6421 dummy_9.n304 dummy_9.n303 0.849769
R6422 dummy_9.n303 dummy_9.n302 0.849769
R6423 dummy_9.n302 dummy_9.n301 0.849769
R6424 dummy_9.n301 dummy_9.n300 0.849769
R6425 dummy_9.n300 dummy_9.n299 0.849769
R6426 dummy_9.n299 dummy_9.n298 0.849769
R6427 dummy_9.n298 dummy_9.n297 0.849769
R6428 dummy_9.n297 dummy_9.n296 0.849769
R6429 dummy_9.n296 dummy_9.n295 0.849769
R6430 dummy_9.n295 dummy_9.n294 0.849769
R6431 dummy_9.n294 dummy_9.n293 0.849769
R6432 dummy_9.n293 dummy_9.n292 0.849769
R6433 dummy_9.n292 dummy_9.n291 0.849769
R6434 dummy_9.n291 dummy_9.n290 0.849769
R6435 dummy_9.n290 dummy_9.n289 0.849769
R6436 dummy_9.n289 dummy_9.n288 0.849769
R6437 dummy_9.n288 dummy_9.n287 0.849769
R6438 dummy_9.n287 dummy_9.n286 0.849769
R6439 dummy_9.n286 dummy_9.n285 0.849769
R6440 dummy_9.n285 dummy_9.n284 0.849769
R6441 dummy_9.n284 dummy_9.n283 0.849769
R6442 dummy_9.n283 dummy_9.n282 0.849769
R6443 dummy_9.n282 dummy_9.n281 0.849769
R6444 dummy_9.n281 dummy_9.n280 0.849769
R6445 dummy_9.n280 dummy_9.n279 0.849769
R6446 dummy_9.n279 dummy_9.n278 0.849769
R6447 dummy_9.n278 dummy_9.n277 0.849769
R6448 dummy_9.n277 dummy_9.n276 0.849769
R6449 dummy_9.n276 dummy_9.n275 0.849769
R6450 dummy_9.n275 dummy_9.n274 0.849769
R6451 dummy_9.n274 dummy_9.n273 0.849769
R6452 dummy_9.n273 dummy_9.n272 0.849769
R6453 dummy_9.n272 dummy_9.n271 0.849769
R6454 dummy_9.n271 dummy_9.n270 0.849769
R6455 dummy_9.n270 dummy_9.n269 0.849769
R6456 dummy_9.n269 dummy_9.n268 0.849769
R6457 dummy_9.n268 dummy_9.n267 0.849769
R6458 dummy_9.n267 dummy_9.n266 0.849769
R6459 dummy_9.n266 dummy_9.n265 0.849769
R6460 dummy_9.n265 dummy_9.n264 0.849769
R6461 dummy_9.n264 dummy_9.n263 0.849769
R6462 dummy_9.n263 dummy_9.n262 0.849769
R6463 dummy_9.n262 dummy_9.n261 0.849769
R6464 dummy_9.n261 dummy_9.n260 0.849769
R6465 dummy_9.n260 dummy_9.n259 0.849769
R6466 dummy_9.n259 dummy_9.n258 0.849769
R6467 dummy_9.n258 dummy_9.n257 0.849769
R6468 dummy_9.n257 dummy_9.n256 0.849769
R6469 dummy_9.n256 dummy_9.n255 0.849769
R6470 dummy_9.n255 dummy_9.n254 0.849769
R6471 dummy_9.n254 dummy_9.n253 0.849769
R6472 dummy_9.n253 dummy_9.n252 0.849769
R6473 dummy_9.n252 dummy_9.n251 0.849769
R6474 dummy_9.n251 dummy_9.n250 0.849769
R6475 dummy_9.n250 dummy_9.n249 0.849769
R6476 dummy_9.n249 dummy_9.n248 0.849769
R6477 dummy_9.n248 dummy_9.n247 0.849769
R6478 dummy_9.n247 dummy_9.n246 0.849769
R6479 dummy_9.n246 dummy_9.n245 0.849769
R6480 dummy_9.n245 dummy_9.n244 0.849769
R6481 dummy_9.n244 dummy_9.n243 0.849769
R6482 dummy_9.n243 dummy_9.n242 0.849769
R6483 dummy_9.n242 dummy_9.n241 0.849769
R6484 dummy_9.n241 dummy_9.n240 0.849769
R6485 dummy_9.n240 dummy_9.n239 0.849769
R6486 dummy_9.n239 dummy_9.n238 0.849769
R6487 dummy_9.n238 dummy_9.n237 0.849769
R6488 dummy_9.n237 dummy_9.n236 0.849769
R6489 dummy_9.n236 dummy_9.n235 0.849769
R6490 dummy_9.n235 dummy_9.n234 0.849769
R6491 dummy_9.n234 dummy_9.n233 0.849769
R6492 dummy_9.n233 dummy_9.n232 0.849769
R6493 dummy_9.n232 dummy_9.n231 0.849769
R6494 dummy_9.n231 dummy_9.n230 0.849769
R6495 dummy_9.n230 dummy_9.n229 0.849769
R6496 dummy_9.n3 dummy_9.n2 0.849769
R6497 dummy_9.n4 dummy_9.n3 0.849769
R6498 dummy_9.n446 dummy_9.n445 0.849769
R6499 dummy_9.n445 dummy_9.n444 0.849769
R6500 dummy_9.n444 dummy_9.n443 0.849769
R6501 dummy_9.n443 dummy_9.n442 0.849769
R6502 dummy_9.n442 dummy_9.n441 0.849769
R6503 dummy_9.n441 dummy_9.n440 0.849769
R6504 dummy_9.n440 dummy_9.n439 0.849769
R6505 dummy_9.n439 dummy_9.n438 0.849769
R6506 dummy_9.n438 dummy_9.n437 0.849769
R6507 dummy_9.n437 dummy_9.n436 0.849769
R6508 dummy_9.n436 dummy_9.n435 0.849769
R6509 dummy_9.n435 dummy_9.n434 0.849769
R6510 dummy_9.n434 dummy_9.n433 0.849769
R6511 dummy_9.n433 dummy_9.n432 0.849769
R6512 dummy_9.n432 dummy_9.n431 0.849769
R6513 dummy_9.n431 dummy_9.n430 0.849769
R6514 dummy_9.n430 dummy_9.n429 0.849769
R6515 dummy_9.n429 dummy_9.n428 0.849769
R6516 dummy_9.n428 dummy_9.n427 0.849769
R6517 dummy_9.n427 dummy_9.n426 0.849769
R6518 dummy_9.n426 dummy_9.n425 0.849769
R6519 dummy_9.n425 dummy_9.n424 0.849769
R6520 dummy_9.n424 dummy_9.n423 0.849769
R6521 dummy_9.n423 dummy_9.n422 0.849769
R6522 dummy_9.n422 dummy_9.n421 0.849769
R6523 dummy_9.n421 dummy_9.n420 0.849769
R6524 dummy_9.n420 dummy_9.n419 0.849769
R6525 dummy_9.n419 dummy_9.n418 0.849769
R6526 dummy_9.n418 dummy_9.n417 0.849769
R6527 dummy_9.n417 dummy_9.n416 0.849769
R6528 dummy_9.n416 dummy_9.n415 0.849769
R6529 dummy_9.n415 dummy_9.n414 0.849769
R6530 dummy_9.n414 dummy_9.n413 0.849769
R6531 dummy_9.n413 dummy_9.n412 0.849769
R6532 dummy_9.n412 dummy_9.n411 0.849769
R6533 dummy_9.n411 dummy_9.n410 0.849769
R6534 dummy_9.n410 dummy_9.n409 0.849769
R6535 dummy_9.n409 dummy_9.n408 0.849769
R6536 dummy_9.n408 dummy_9.n407 0.849769
R6537 dummy_9.n407 dummy_9.n406 0.849769
R6538 dummy_9.n406 dummy_9.n405 0.849769
R6539 dummy_9.n405 dummy_9.n404 0.849769
R6540 dummy_9.n404 dummy_9.n403 0.849769
R6541 dummy_9.n403 dummy_9.n402 0.849769
R6542 dummy_9.n402 dummy_9.n401 0.849769
R6543 dummy_9.n401 dummy_9.n400 0.849769
R6544 dummy_9.n400 dummy_9.n399 0.849769
R6545 dummy_9.n399 dummy_9.n398 0.849769
R6546 dummy_9.n398 dummy_9.n397 0.849769
R6547 dummy_9.n397 dummy_9.n396 0.849769
R6548 dummy_9.n396 dummy_9.n395 0.849769
R6549 dummy_9.n395 dummy_9.n394 0.849769
R6550 dummy_9.n394 dummy_9.n393 0.849769
R6551 dummy_9.n393 dummy_9.n392 0.849769
R6552 dummy_9.n392 dummy_9.n391 0.849769
R6553 dummy_9.n391 dummy_9.n390 0.849769
R6554 dummy_9.n390 dummy_9.n389 0.849769
R6555 dummy_9.n389 dummy_9.n388 0.849769
R6556 dummy_9.n388 dummy_9.n387 0.849769
R6557 dummy_9.n387 dummy_9.n386 0.849769
R6558 dummy_9.n386 dummy_9.n385 0.849769
R6559 dummy_9.n385 dummy_9.n384 0.849769
R6560 dummy_9.n384 dummy_9.n383 0.849769
R6561 dummy_9.n383 dummy_9.n382 0.849769
R6562 dummy_9.n382 dummy_9.n381 0.849769
R6563 dummy_9.n381 dummy_9.n380 0.849769
R6564 dummy_9.n380 dummy_9.n379 0.849769
R6565 dummy_9.n379 dummy_9.n378 0.849769
R6566 dummy_9.n378 dummy_9.n377 0.849769
R6567 dummy_9.n377 dummy_9.n376 0.849769
R6568 dummy_9.n376 dummy_9.n375 0.849769
R6569 dummy_9.n375 dummy_9.n374 0.849769
R6570 dummy_9.n374 dummy_9.n373 0.849769
R6571 dummy_9.n373 dummy_9.n372 0.849769
R6572 dummy_9.n372 dummy_9.n371 0.849769
R6573 dummy_9.n5 dummy_9.n4 0.838728
R6574 dummy_9.n25 dummy_9.n24 0.789389
R6575 dummy_9.n26 dummy_9.n25 0.789389
R6576 dummy_9.n27 dummy_9.n26 0.789389
R6577 dummy_9.n28 dummy_9.n27 0.789389
R6578 dummy_9.n29 dummy_9.n28 0.789389
R6579 dummy_9.n30 dummy_9.n29 0.789389
R6580 dummy_9.n31 dummy_9.n30 0.789389
R6581 dummy_9.n32 dummy_9.n31 0.789389
R6582 dummy_9.n33 dummy_9.n32 0.789389
R6583 dummy_9.n34 dummy_9.n33 0.789389
R6584 dummy_9.n35 dummy_9.n34 0.789389
R6585 dummy_9.n36 dummy_9.n35 0.789389
R6586 dummy_9.n37 dummy_9.n36 0.789389
R6587 dummy_9.n38 dummy_9.n37 0.789389
R6588 dummy_9.n39 dummy_9.n38 0.789389
R6589 dummy_9.n40 dummy_9.n39 0.789389
R6590 dummy_9.n41 dummy_9.n40 0.789389
R6591 dummy_9.n42 dummy_9.n41 0.789389
R6592 dummy_9.n43 dummy_9.n42 0.789389
R6593 dummy_9.n44 dummy_9.n43 0.789389
R6594 dummy_9.n45 dummy_9.n44 0.789389
R6595 dummy_9.n46 dummy_9.n45 0.789389
R6596 dummy_9.n47 dummy_9.n46 0.789389
R6597 dummy_9.n48 dummy_9.n47 0.789389
R6598 dummy_9.n49 dummy_9.n48 0.789389
R6599 dummy_9.n50 dummy_9.n49 0.789389
R6600 dummy_9.n51 dummy_9.n50 0.789389
R6601 dummy_9.n52 dummy_9.n51 0.789389
R6602 dummy_9.n53 dummy_9.n52 0.789389
R6603 dummy_9.n54 dummy_9.n53 0.789389
R6604 dummy_9.n55 dummy_9.n54 0.789389
R6605 dummy_9.n56 dummy_9.n55 0.789389
R6606 dummy_9.n57 dummy_9.n56 0.789389
R6607 dummy_9.n58 dummy_9.n57 0.789389
R6608 dummy_9.n59 dummy_9.n58 0.789389
R6609 dummy_9.n60 dummy_9.n59 0.789389
R6610 dummy_9.n61 dummy_9.n60 0.789389
R6611 dummy_9.n62 dummy_9.n61 0.789389
R6612 dummy_9.n63 dummy_9.n62 0.789389
R6613 dummy_9.n64 dummy_9.n63 0.789389
R6614 dummy_9.n65 dummy_9.n64 0.789389
R6615 dummy_9.n66 dummy_9.n65 0.789389
R6616 dummy_9.n67 dummy_9.n66 0.789389
R6617 dummy_9.n68 dummy_9.n67 0.789389
R6618 dummy_9.n69 dummy_9.n68 0.789389
R6619 dummy_9.n70 dummy_9.n69 0.789389
R6620 dummy_9.n71 dummy_9.n70 0.789389
R6621 dummy_9.n72 dummy_9.n71 0.789389
R6622 dummy_9.n73 dummy_9.n72 0.789389
R6623 dummy_9.n74 dummy_9.n73 0.789389
R6624 dummy_9.n75 dummy_9.n74 0.789389
R6625 dummy_9.n76 dummy_9.n75 0.789389
R6626 dummy_9.n77 dummy_9.n76 0.789389
R6627 dummy_9.n78 dummy_9.n77 0.789389
R6628 dummy_9.n79 dummy_9.n78 0.789389
R6629 dummy_9.n80 dummy_9.n79 0.789389
R6630 dummy_9.n81 dummy_9.n80 0.789389
R6631 dummy_9.n82 dummy_9.n81 0.789389
R6632 dummy_9.n83 dummy_9.n82 0.789389
R6633 dummy_9.n84 dummy_9.n83 0.789389
R6634 dummy_9.n85 dummy_9.n84 0.789389
R6635 dummy_9.n86 dummy_9.n85 0.789389
R6636 dummy_9.n87 dummy_9.n86 0.789389
R6637 dummy_9.n88 dummy_9.n87 0.789389
R6638 dummy_9.n89 dummy_9.n88 0.789389
R6639 dummy_9.n90 dummy_9.n89 0.789389
R6640 dummy_9.n91 dummy_9.n90 0.789389
R6641 dummy_9.n92 dummy_9.n91 0.789389
R6642 dummy_9.n93 dummy_9.n92 0.789389
R6643 dummy_9.n94 dummy_9.n93 0.789389
R6644 dummy_9.n95 dummy_9.n94 0.789389
R6645 dummy_9.n96 dummy_9.n95 0.789389
R6646 dummy_9.n97 dummy_9.n96 0.789389
R6647 dummy_9.n98 dummy_9.n97 0.789389
R6648 dummy_9.n99 dummy_9.n98 0.789389
R6649 dummy_9.n100 dummy_9.n99 0.789389
R6650 dummy_9.n101 dummy_9.n100 0.789389
R6651 dummy_9.n102 dummy_9.n101 0.789389
R6652 dummy_9.n103 dummy_9.n102 0.789389
R6653 dummy_9.n104 dummy_9.n103 0.789389
R6654 dummy_9.n130 dummy_9.n129 0.789389
R6655 dummy_9.n131 dummy_9.n130 0.789389
R6656 dummy_9.n132 dummy_9.n131 0.789389
R6657 dummy_9.n133 dummy_9.n132 0.789389
R6658 dummy_9.n134 dummy_9.n133 0.789389
R6659 dummy_9.n135 dummy_9.n134 0.789389
R6660 dummy_9.n136 dummy_9.n135 0.789389
R6661 dummy_9.n137 dummy_9.n136 0.789389
R6662 dummy_9.n138 dummy_9.n137 0.789389
R6663 dummy_9.n139 dummy_9.n138 0.789389
R6664 dummy_9.n140 dummy_9.n139 0.789389
R6665 dummy_9.n141 dummy_9.n140 0.789389
R6666 dummy_9.n142 dummy_9.n141 0.789389
R6667 dummy_9.n143 dummy_9.n142 0.789389
R6668 dummy_9.n144 dummy_9.n143 0.789389
R6669 dummy_9.n145 dummy_9.n144 0.789389
R6670 dummy_9.n146 dummy_9.n145 0.789389
R6671 dummy_9.n147 dummy_9.n146 0.789389
R6672 dummy_9.n148 dummy_9.n147 0.789389
R6673 dummy_9.n149 dummy_9.n148 0.789389
R6674 dummy_9.n150 dummy_9.n149 0.789389
R6675 dummy_9.n151 dummy_9.n150 0.789389
R6676 dummy_9.n152 dummy_9.n151 0.789389
R6677 dummy_9.n153 dummy_9.n152 0.789389
R6678 dummy_9.n154 dummy_9.n153 0.789389
R6679 dummy_9.n155 dummy_9.n154 0.789389
R6680 dummy_9.n156 dummy_9.n155 0.789389
R6681 dummy_9.n157 dummy_9.n156 0.789389
R6682 dummy_9.n158 dummy_9.n157 0.789389
R6683 dummy_9.n159 dummy_9.n158 0.789389
R6684 dummy_9.n160 dummy_9.n159 0.789389
R6685 dummy_9.n161 dummy_9.n160 0.789389
R6686 dummy_9.n162 dummy_9.n161 0.789389
R6687 dummy_9.n163 dummy_9.n162 0.789389
R6688 dummy_9.n164 dummy_9.n163 0.789389
R6689 dummy_9.n165 dummy_9.n164 0.789389
R6690 dummy_9.n166 dummy_9.n165 0.789389
R6691 dummy_9.n167 dummy_9.n166 0.789389
R6692 dummy_9.n168 dummy_9.n167 0.789389
R6693 dummy_9.n169 dummy_9.n168 0.789389
R6694 dummy_9.n170 dummy_9.n169 0.789389
R6695 dummy_9.n171 dummy_9.n170 0.789389
R6696 dummy_9.n172 dummy_9.n171 0.789389
R6697 dummy_9.n173 dummy_9.n172 0.789389
R6698 dummy_9.n174 dummy_9.n173 0.789389
R6699 dummy_9.n175 dummy_9.n174 0.789389
R6700 dummy_9.n176 dummy_9.n175 0.789389
R6701 dummy_9.n177 dummy_9.n176 0.789389
R6702 dummy_9.n178 dummy_9.n177 0.789389
R6703 dummy_9.n179 dummy_9.n178 0.789389
R6704 dummy_9.n180 dummy_9.n179 0.789389
R6705 dummy_9.n181 dummy_9.n180 0.789389
R6706 dummy_9.n182 dummy_9.n181 0.789389
R6707 dummy_9.n183 dummy_9.n182 0.789389
R6708 dummy_9.n184 dummy_9.n183 0.789389
R6709 dummy_9.n185 dummy_9.n184 0.789389
R6710 dummy_9.n186 dummy_9.n185 0.789389
R6711 dummy_9.n187 dummy_9.n186 0.789389
R6712 dummy_9.n188 dummy_9.n187 0.789389
R6713 dummy_9.n189 dummy_9.n188 0.789389
R6714 dummy_9.n190 dummy_9.n189 0.789389
R6715 dummy_9.n191 dummy_9.n190 0.789389
R6716 dummy_9.n192 dummy_9.n191 0.789389
R6717 dummy_9.n193 dummy_9.n192 0.789389
R6718 dummy_9.n194 dummy_9.n193 0.789389
R6719 dummy_9.n195 dummy_9.n194 0.789389
R6720 dummy_9.n196 dummy_9.n195 0.789389
R6721 dummy_9.n197 dummy_9.n196 0.789389
R6722 dummy_9.n198 dummy_9.n197 0.789389
R6723 dummy_9.n199 dummy_9.n198 0.789389
R6724 dummy_9.n200 dummy_9.n199 0.789389
R6725 dummy_9.n201 dummy_9.n200 0.789389
R6726 dummy_9.n202 dummy_9.n201 0.789389
R6727 dummy_9.n203 dummy_9.n202 0.789389
R6728 dummy_9.n204 dummy_9.n203 0.789389
R6729 dummy_9.n205 dummy_9.n204 0.789389
R6730 dummy_9.n206 dummy_9.n205 0.789389
R6731 dummy_9.n207 dummy_9.n206 0.789389
R6732 dummy_9.n208 dummy_9.n207 0.789389
R6733 dummy_9.n209 dummy_9.n208 0.789389
R6734 dummy_9.n210 dummy_9.n209 0.789389
R6735 dummy_9.n211 dummy_9.n210 0.789389
R6736 dummy_9.n212 dummy_9.n211 0.789389
R6737 dummy_9.n213 dummy_9.n212 0.789389
R6738 dummy_9.n214 dummy_9.n213 0.789389
R6739 dummy_9.n215 dummy_9.n214 0.789389
R6740 dummy_9.n216 dummy_9.n215 0.789389
R6741 dummy_9.n217 dummy_9.n216 0.789389
R6742 dummy_9.n218 dummy_9.n217 0.789389
R6743 dummy_9.n219 dummy_9.n218 0.789389
R6744 dummy_9.n220 dummy_9.n219 0.789389
R6745 dummy_9.n221 dummy_9.n220 0.789389
R6746 dummy_9.n222 dummy_9.n221 0.789389
R6747 dummy_9.n223 dummy_9.n222 0.789389
R6748 dummy_9.n224 dummy_9.n223 0.789389
R6749 dummy_9.n225 dummy_9.n224 0.789389
R6750 dummy_9.n226 dummy_9.n225 0.789389
R6751 dummy_9.n227 dummy_9.n226 0.789389
R6752 dummy_9.n228 dummy_9.n227 0.789389
R6753 dummy_9.n105 dummy_9.n104 0.779191
R6754 dummy_9.n129 dummy_9.n128 0.779188
R6755 dummy_9.n326 dummy_9.n325 0.750892
R6756 dummy_9.n7 dummy_9.n6 0.740222
R6757 dummy_9.n11 dummy_9.n10 0.740222
R6758 dummy_9.n13 dummy_9.n12 0.740222
R6759 dummy_9.n19 dummy_9.n18 0.740222
R6760 dummy_9.n20 dummy_9.n19 0.735222
R6761 dummy_9.n24 dummy_9.n23 0.723556
R6762 dummy_9.n21 dummy_9.n20 0.703556
R6763 dummy_9.n8 dummy_9.n7 0.698556
R6764 dummy_9.n9 dummy_9.n8 0.698556
R6765 dummy_9.n10 dummy_9.n9 0.698556
R6766 dummy_9.n22 dummy_9.n21 0.698556
R6767 dummy_9.n23 dummy_9.n22 0.698556
R6768 dummy_9.n14 dummy_9.n13 0.698556
R6769 dummy_9.n15 dummy_9.n14 0.698556
R6770 dummy_9.n16 dummy_9.n15 0.698556
R6771 dummy_9.n17 dummy_9.n16 0.698556
R6772 dummy_9.n18 dummy_9.n17 0.698556
R6773 dummy_9.n12 dummy_9.n11 0.656889
R6774 dummy_9.n346 dummy_9.n345 0.464029
R6775 dummy_9.n344 dummy_9.n343 0.464029
R6776 dummy_9.n342 dummy_9.n341 0.464029
R6777 dummy_9.n340 dummy_9.n339 0.464029
R6778 dummy_9.n338 dummy_9.n337 0.464029
R6779 dummy_9.n336 dummy_9.n335 0.464029
R6780 dummy_9.n334 dummy_9.n333 0.464029
R6781 dummy_9.n332 dummy_9.n331 0.464029
R6782 dummy_9.n330 dummy_9.n329 0.464029
R6783 dummy_9.n328 dummy_9.n327 0.464029
R6784 dummy_9.n127 dummy_9.n126 0.464029
R6785 dummy_9.n125 dummy_9.n124 0.464029
R6786 dummy_9.n123 dummy_9.n122 0.464029
R6787 dummy_9.n121 dummy_9.n120 0.464029
R6788 dummy_9.n119 dummy_9.n118 0.464029
R6789 dummy_9.n117 dummy_9.n116 0.464029
R6790 dummy_9.n115 dummy_9.n114 0.464029
R6791 dummy_9.n113 dummy_9.n112 0.464029
R6792 dummy_9.n111 dummy_9.n110 0.464029
R6793 dummy_9.n109 dummy_9.n108 0.464029
R6794 dummy_9.n107 dummy_9.n106 0.464029
R6795 dummy_9 dummy_9.n228 0.449111
R6796 dummy_9.n1 dummy_9.n347 0.343416
R6797 dummy_9 dummy_9.n447 0.248168
R6798 dummy_9.n0 dummy_9.n1 0.0510086
R6799 dummy_9.n106 dummy_9.n105 0.02299
R6800 bias3.n8 bias3.t42 65.7904
R6801 bias3.n9 bias3.t46 43.8281
R6802 bias3.n30 bias3.t44 43.3905
R6803 bias3.n35 bias3.t47 43.3905
R6804 bias3.n27 bias3.t57 43.3864
R6805 bias3.n25 bias3.t43 43.3864
R6806 bias3.n17 bias3.t56 43.3861
R6807 bias3.n16 bias3.t49 43.3861
R6808 bias3.n15 bias3.t55 43.3861
R6809 bias3.n28 bias3.t54 43.3861
R6810 bias3.n26 bias3.t41 43.3861
R6811 bias3.n14 bias3.t45 43.3861
R6812 bias3.n13 bias3.t48 43.3847
R6813 bias3 bias3.n52 37.6626
R6814 bias3.n1 bias3.t4 22.674
R6815 bias3.n9 bias3.t40 21.5536
R6816 bias3.n10 bias3.t53 21.5536
R6817 bias3.n11 bias3.t51 21.5536
R6818 bias3.n12 bias3.t38 21.5536
R6819 bias3.n34 bias3.t58 21.5536
R6820 bias3.n33 bias3.t50 21.5536
R6821 bias3.n32 bias3.t52 21.5536
R6822 bias3.n31 bias3.t39 21.5536
R6823 bias3.n3 bias3.t6 21.4458
R6824 bias3.n2 bias3.t0 21.4435
R6825 bias3.n1 bias3.t2 21.4435
R6826 bias3.n37 bias3.n36 16.2841
R6827 bias3.n4 bias3.t5 15.1153
R6828 bias3.n6 bias3.t7 13.9238
R6829 bias3.n5 bias3.t1 13.9238
R6830 bias3.n4 bias3.t3 13.9238
R6831 bias3.n50 bias3.t28 6.90631
R6832 bias3.n50 bias3.t36 6.90131
R6833 bias3.n41 bias3.t12 6.84109
R6834 bias3.n41 bias3.t17 6.83609
R6835 bias3.n52 bias3.t29 6.83022
R6836 bias3.n52 bias3.t15 6.82522
R6837 bias3.n38 bias3.t20 6.81935
R6838 bias3.n38 bias3.t19 6.81435
R6839 bias3.n49 bias3.t37 6.80848
R6840 bias3.n49 bias3.t33 6.80348
R6841 bias3.n46 bias3.t27 6.78674
R6842 bias3.n46 bias3.t35 6.78174
R6843 bias3.n43 bias3.t32 6.76501
R6844 bias3.n43 bias3.t24 6.76001
R6845 bias3.n40 bias3.t13 6.74327
R6846 bias3.n40 bias3.t18 6.73827
R6847 bias3.n51 bias3.t16 6.7324
R6848 bias3.n51 bias3.t9 6.7274
R6849 bias3.n48 bias3.t14 6.71066
R6850 bias3.n48 bias3.t8 6.70566
R6851 bias3.n45 bias3.t11 6.68892
R6852 bias3.n45 bias3.t23 6.68392
R6853 bias3.n42 bias3.t31 6.66718
R6854 bias3.n42 bias3.t34 6.66218
R6855 bias3.n39 bias3.t10 6.64544
R6856 bias3.n39 bias3.t22 6.64044
R6857 bias3.n47 bias3.t25 6.61283
R6858 bias3.n47 bias3.t26 6.60783
R6859 bias3.n44 bias3.t30 6.59109
R6860 bias3.n44 bias3.t21 6.58609
R6861 bias3.n37 bias3.n8 4.44926
R6862 bias3.n8 bias3.n7 2.93009
R6863 bias3.n2 bias3.n1 1.231
R6864 bias3.n3 bias3.n2 1.22634
R6865 bias3.n5 bias3.n4 1.19203
R6866 bias3.n6 bias3.n5 1.19203
R6867 bias3.n7 bias3.n3 0.890317
R6868 bias3.n51 bias3.n50 0.739136
R6869 bias3.n47 bias3.n46 0.739136
R6870 bias3.n44 bias3.n43 0.739136
R6871 bias3.n42 bias3.n41 0.739136
R6872 bias3.n39 bias3.n38 0.739136
R6873 bias3.n10 bias3.n9 0.729127
R6874 bias3.n11 bias3.n10 0.729127
R6875 bias3.n12 bias3.n11 0.729127
R6876 bias3.n34 bias3.n33 0.729127
R6877 bias3.n33 bias3.n32 0.729127
R6878 bias3.n32 bias3.n31 0.729127
R6879 bias3.n14 bias3.n13 0.696048
R6880 bias3.n20 bias3.n19 0.692795
R6881 bias3.n27 bias3.n26 0.692795
R6882 bias3.n21 bias3.n20 0.692544
R6883 bias3.n22 bias3.n21 0.692544
R6884 bias3.n15 bias3.n14 0.692338
R6885 bias3.n16 bias3.n15 0.692338
R6886 bias3.n17 bias3.n16 0.692338
R6887 bias3.n26 bias3.n25 0.692086
R6888 bias3.n28 bias3.n27 0.692086
R6889 bias3.n36 bias3.n17 0.689439
R6890 bias3.n52 bias3.n51 0.682318
R6891 bias3.n50 bias3.n49 0.682318
R6892 bias3.n49 bias3.n48 0.682318
R6893 bias3.n48 bias3.n47 0.682318
R6894 bias3.n46 bias3.n45 0.682318
R6895 bias3.n45 bias3.n44 0.682318
R6896 bias3.n43 bias3.n42 0.682318
R6897 bias3.n41 bias3.n40 0.682318
R6898 bias3.n40 bias3.n39 0.682318
R6899 bias3.n13 bias3.n12 1.01342
R6900 bias3.n35 bias3.n0 0.567567
R6901 bias3.n25 bias3.n24 0.56039
R6902 bias3.n19 bias3.n18 0.559932
R6903 bias3.n29 bias3.n28 0.558947
R6904 bias3.n23 bias3.n22 0.558696
R6905 bias3.n7 bias3.n6 0.418141
R6906 bias3.n0 bias3.n34 0.410126
R6907 bias3.n30 bias3.n29 0.134875
R6908 bias3 bias3.n37 0.128769
R6909 bias3.n36 bias3.n35 0.00280782
R6910 bias3.n31 bias3.n30 0.439043
R6911 bias3.n0 bias3.n23 0.170257
R6912 dummy_4.n19 dummy_4.t19 13.9463
R6913 dummy_4.n21 dummy_4.t7 13.9463
R6914 dummy_4.n20 dummy_4.t18 13.9459
R6915 dummy_4.n22 dummy_4.t6 13.9459
R6916 dummy_4.n17 dummy_4.t5 13.933
R6917 dummy_4.n28 dummy_4.t8 13.932
R6918 dummy_4.n30 dummy_4.t2 13.932
R6919 dummy_4.n32 dummy_4.t32 13.932
R6920 dummy_4.n34 dummy_4.t30 13.932
R6921 dummy_4.n18 dummy_4.t4 13.932
R6922 dummy_4.n24 dummy_4.t26 13.932
R6923 dummy_4.n27 dummy_4.t9 13.9319
R6924 dummy_4.n29 dummy_4.t3 13.9319
R6925 dummy_4.n31 dummy_4.t33 13.9319
R6926 dummy_4.n33 dummy_4.t31 13.9319
R6927 dummy_4.n23 dummy_4.t27 13.9319
R6928 dummy_4.n2 dummy_4.t22 13.9315
R6929 dummy_4.n16 dummy_4.t23 13.931
R6930 dummy_4.n3 dummy_4.t21 13.9305
R6931 dummy_4.n25 dummy_4.t20 13.9305
R6932 dummy_4.n35 dummy_4.t24 13.9259
R6933 dummy_4.n1 dummy_4.t28 13.9259
R6934 dummy_4.n0 dummy_4.t25 13.9259
R6935 dummy_4.n26 dummy_4.t29 13.9258
R6936 dummy_4.n6 dummy_4.t15 13.9238
R6937 dummy_4.n5 dummy_4.t11 13.9238
R6938 dummy_4.n4 dummy_4.t35 13.9238
R6939 dummy_4.n8 dummy_4.t36 13.9238
R6940 dummy_4.n9 dummy_4.t12 13.9238
R6941 dummy_4.n10 dummy_4.t16 13.9238
R6942 dummy_4.n11 dummy_4.t0 13.9238
R6943 dummy_4.n15 dummy_4.t1 13.9238
R6944 dummy_4.n14 dummy_4.t17 13.9238
R6945 dummy_4.n13 dummy_4.t13 13.9238
R6946 dummy_4.n12 dummy_4.t37 13.9238
R6947 dummy_4.n39 dummy_4.t38 13.9238
R6948 dummy_4.n38 dummy_4.t14 13.9238
R6949 dummy_4.n37 dummy_4.t10 13.9238
R6950 dummy_4.n36 dummy_4.t34 13.9238
R6951 dummy_4.n7 dummy_4.t39 13.9238
R6952 dummy_4.n13 dummy_4.n12 1.50979
R6953 dummy_4.n14 dummy_4.n13 1.50979
R6954 dummy_4.n15 dummy_4.n14 1.50979
R6955 dummy_4.n5 dummy_4.n4 1.50979
R6956 dummy_4.n6 dummy_4.n5 1.50979
R6957 dummy_4.n7 dummy_4.n6 1.50979
R6958 dummy_4.n37 dummy_4.n36 1.46687
R6959 dummy_4.n38 dummy_4.n37 1.46687
R6960 dummy_4.n39 dummy_4.n38 1.46687
R6961 dummy_4.n11 dummy_4.n10 1.46687
R6962 dummy_4.n10 dummy_4.n9 1.46687
R6963 dummy_4.n9 dummy_4.n8 1.46687
R6964 dummy_4.n16 dummy_4.n15 1.46027
R6965 dummy_4.n3 dummy_4.n7 1.45167
R6966 dummy_4.n36 dummy_4.n35 1.42112
R6967 dummy_4.n2 dummy_4.n11 1.41789
R6968 dummy_4 dummy_4.n39 0.821185
R6969 dummy_4 dummy_4.n25 0.597208
R6970 dummy_4.n2 dummy_4.n16 0.481643
R6971 dummy_4.n18 dummy_4.n17 0.434926
R6972 dummy_4.n25 dummy_4.n3 0.410477
R6973 dummy_4.n22 dummy_4.n21 0.388284
R6974 dummy_4.n20 dummy_4.n19 0.388284
R6975 dummy_4.n24 dummy_4.n23 0.366986
R6976 dummy_4.n1 dummy_4.n26 0.308718
R6977 dummy_4.n17 dummy_4.n2 0.296602
R6978 dummy_4.n23 dummy_4.n22 0.283532
R6979 dummy_4.n35 dummy_4.n0 0.268628
R6980 dummy_4.n34 dummy_4.n33 0.264861
R6981 dummy_4.n32 dummy_4.n31 0.264861
R6982 dummy_4.n30 dummy_4.n29 0.264861
R6983 dummy_4.n28 dummy_4.n27 0.264861
R6984 dummy_4.n3 dummy_4.n24 0.250346
R6985 dummy_4.n21 dummy_4.n20 0.249454
R6986 dummy_4.n19 dummy_4.n18 0.249454
R6987 dummy_4.n27 dummy_4.n1 0.220446
R6988 dummy_4.n0 dummy_4.n34 0.22044
R6989 dummy_4.n33 dummy_4.n32 0.214688
R6990 dummy_4.n31 dummy_4.n30 0.214688
R6991 dummy_4.n29 dummy_4.n28 0.214688
R6992 VB_A.n67 VB_A.t16 13.7936
R6993 VB_A.n50 VB_A.t75 13.7936
R6994 VB_A.n33 VB_A.t36 13.7936
R6995 VB_A.n16 VB_A.t89 13.7936
R6996 VB_A.n84 VB_A.t64 13.7927
R6997 VB_A.n0 VB_A.t93 13.7927
R6998 VB_A.n84 VB_A.t12 13.5352
R6999 VB_A.n85 VB_A.t88 13.5352
R7000 VB_A.n86 VB_A.t67 13.5352
R7001 VB_A.n87 VB_A.t43 13.5352
R7002 VB_A.n88 VB_A.t21 13.5352
R7003 VB_A.n89 VB_A.t41 13.5352
R7004 VB_A.n90 VB_A.t24 13.5352
R7005 VB_A.n91 VB_A.t71 13.5352
R7006 VB_A.n92 VB_A.t23 13.5352
R7007 VB_A.n93 VB_A.t100 13.5352
R7008 VB_A.n94 VB_A.t4 13.5352
R7009 VB_A.n95 VB_A.t54 13.5352
R7010 VB_A.n96 VB_A.t1 13.5352
R7011 VB_A.n97 VB_A.t53 13.5352
R7012 VB_A.n98 VB_A.t35 13.5352
R7013 VB_A.n99 VB_A.t81 13.5352
R7014 VB_A.n67 VB_A.t26 13.5352
R7015 VB_A.n68 VB_A.t74 13.5352
R7016 VB_A.n69 VB_A.t85 13.5352
R7017 VB_A.n70 VB_A.t29 13.5352
R7018 VB_A.n71 VB_A.t5 13.5352
R7019 VB_A.n72 VB_A.t58 13.5352
R7020 VB_A.n73 VB_A.t11 13.5352
R7021 VB_A.n74 VB_A.t87 13.5352
R7022 VB_A.n75 VB_A.t8 13.5352
R7023 VB_A.n76 VB_A.t86 13.5352
R7024 VB_A.n77 VB_A.t96 13.5352
R7025 VB_A.n78 VB_A.t40 13.5352
R7026 VB_A.n79 VB_A.t17 13.5352
R7027 VB_A.n80 VB_A.t38 13.5352
R7028 VB_A.n81 VB_A.t22 13.5352
R7029 VB_A.n82 VB_A.t99 13.5352
R7030 VB_A.n50 VB_A.t90 13.5352
R7031 VB_A.n51 VB_A.t34 13.5352
R7032 VB_A.n52 VB_A.t44 13.5352
R7033 VB_A.n53 VB_A.t92 13.5352
R7034 VB_A.n54 VB_A.t65 13.5352
R7035 VB_A.n55 VB_A.t19 13.5352
R7036 VB_A.n56 VB_A.t72 13.5352
R7037 VB_A.n57 VB_A.t47 13.5352
R7038 VB_A.n58 VB_A.t68 13.5352
R7039 VB_A.n59 VB_A.t46 13.5352
R7040 VB_A.n60 VB_A.t56 13.5352
R7041 VB_A.n61 VB_A.t3 13.5352
R7042 VB_A.n62 VB_A.t77 13.5352
R7043 VB_A.n63 VB_A.t0 13.5352
R7044 VB_A.n64 VB_A.t83 13.5352
R7045 VB_A.n65 VB_A.t60 13.5352
R7046 VB_A.n33 VB_A.t49 13.5352
R7047 VB_A.n34 VB_A.t97 13.5352
R7048 VB_A.n35 VB_A.t6 13.5352
R7049 VB_A.n36 VB_A.t52 13.5352
R7050 VB_A.n37 VB_A.t27 13.5352
R7051 VB_A.n38 VB_A.t78 13.5352
R7052 VB_A.n39 VB_A.t33 13.5352
R7053 VB_A.n40 VB_A.t9 13.5352
R7054 VB_A.n41 VB_A.t31 13.5352
R7055 VB_A.n42 VB_A.t7 13.5352
R7056 VB_A.n43 VB_A.t18 13.5352
R7057 VB_A.n44 VB_A.t63 13.5352
R7058 VB_A.n45 VB_A.t39 13.5352
R7059 VB_A.n46 VB_A.t62 13.5352
R7060 VB_A.n47 VB_A.t42 13.5352
R7061 VB_A.n48 VB_A.t20 13.5352
R7062 VB_A.n16 VB_A.t101 13.5352
R7063 VB_A.n17 VB_A.t45 13.5352
R7064 VB_A.n18 VB_A.t55 13.5352
R7065 VB_A.n19 VB_A.t2 13.5352
R7066 VB_A.n20 VB_A.t76 13.5352
R7067 VB_A.n21 VB_A.t32 13.5352
R7068 VB_A.n22 VB_A.t82 13.5352
R7069 VB_A.n23 VB_A.t59 13.5352
R7070 VB_A.n24 VB_A.t79 13.5352
R7071 VB_A.n25 VB_A.t57 13.5352
R7072 VB_A.n26 VB_A.t66 13.5352
R7073 VB_A.n27 VB_A.t15 13.5352
R7074 VB_A.n28 VB_A.t91 13.5352
R7075 VB_A.n29 VB_A.t13 13.5352
R7076 VB_A.n30 VB_A.t94 13.5352
R7077 VB_A.n31 VB_A.t70 13.5352
R7078 VB_A.n0 VB_A.t37 13.5352
R7079 VB_A.n1 VB_A.t14 13.5352
R7080 VB_A.n2 VB_A.t95 13.5352
R7081 VB_A.n3 VB_A.t73 13.5352
R7082 VB_A.n4 VB_A.t48 13.5352
R7083 VB_A.n5 VB_A.t69 13.5352
R7084 VB_A.n6 VB_A.t51 13.5352
R7085 VB_A.n7 VB_A.t98 13.5352
R7086 VB_A.n8 VB_A.t50 13.5352
R7087 VB_A.n9 VB_A.t25 13.5352
R7088 VB_A.n10 VB_A.t30 13.5352
R7089 VB_A.n11 VB_A.t84 13.5352
R7090 VB_A.n12 VB_A.t28 13.5352
R7091 VB_A.n13 VB_A.t80 13.5352
R7092 VB_A.n14 VB_A.t61 13.5352
R7093 VB_A.n15 VB_A.t10 13.5352
R7094 VB_A VB_A.n100 2.25671
R7095 VB_A.n32 VB_A.n15 0.621566
R7096 VB_A.n49 VB_A.n32 0.429071
R7097 VB_A.n66 VB_A.n49 0.429071
R7098 VB_A.n83 VB_A.n66 0.429071
R7099 VB_A.n100 VB_A.n83 0.429071
R7100 VB_A.n85 VB_A.n84 0.257989
R7101 VB_A.n86 VB_A.n85 0.257989
R7102 VB_A.n87 VB_A.n86 0.257989
R7103 VB_A.n88 VB_A.n87 0.257989
R7104 VB_A.n89 VB_A.n88 0.257989
R7105 VB_A.n90 VB_A.n89 0.257989
R7106 VB_A.n91 VB_A.n90 0.257989
R7107 VB_A.n92 VB_A.n91 0.257989
R7108 VB_A.n93 VB_A.n92 0.257989
R7109 VB_A.n94 VB_A.n93 0.257989
R7110 VB_A.n95 VB_A.n94 0.257989
R7111 VB_A.n96 VB_A.n95 0.257989
R7112 VB_A.n97 VB_A.n96 0.257989
R7113 VB_A.n98 VB_A.n97 0.257989
R7114 VB_A.n99 VB_A.n98 0.257989
R7115 VB_A.n68 VB_A.n67 0.257989
R7116 VB_A.n69 VB_A.n68 0.257989
R7117 VB_A.n70 VB_A.n69 0.257989
R7118 VB_A.n71 VB_A.n70 0.257989
R7119 VB_A.n72 VB_A.n71 0.257989
R7120 VB_A.n73 VB_A.n72 0.257989
R7121 VB_A.n74 VB_A.n73 0.257989
R7122 VB_A.n75 VB_A.n74 0.257989
R7123 VB_A.n76 VB_A.n75 0.257989
R7124 VB_A.n77 VB_A.n76 0.257989
R7125 VB_A.n78 VB_A.n77 0.257989
R7126 VB_A.n79 VB_A.n78 0.257989
R7127 VB_A.n80 VB_A.n79 0.257989
R7128 VB_A.n81 VB_A.n80 0.257989
R7129 VB_A.n82 VB_A.n81 0.257989
R7130 VB_A.n51 VB_A.n50 0.257989
R7131 VB_A.n52 VB_A.n51 0.257989
R7132 VB_A.n53 VB_A.n52 0.257989
R7133 VB_A.n54 VB_A.n53 0.257989
R7134 VB_A.n55 VB_A.n54 0.257989
R7135 VB_A.n56 VB_A.n55 0.257989
R7136 VB_A.n57 VB_A.n56 0.257989
R7137 VB_A.n58 VB_A.n57 0.257989
R7138 VB_A.n59 VB_A.n58 0.257989
R7139 VB_A.n60 VB_A.n59 0.257989
R7140 VB_A.n61 VB_A.n60 0.257989
R7141 VB_A.n62 VB_A.n61 0.257989
R7142 VB_A.n63 VB_A.n62 0.257989
R7143 VB_A.n64 VB_A.n63 0.257989
R7144 VB_A.n65 VB_A.n64 0.257989
R7145 VB_A.n34 VB_A.n33 0.257989
R7146 VB_A.n35 VB_A.n34 0.257989
R7147 VB_A.n36 VB_A.n35 0.257989
R7148 VB_A.n37 VB_A.n36 0.257989
R7149 VB_A.n38 VB_A.n37 0.257989
R7150 VB_A.n39 VB_A.n38 0.257989
R7151 VB_A.n40 VB_A.n39 0.257989
R7152 VB_A.n41 VB_A.n40 0.257989
R7153 VB_A.n42 VB_A.n41 0.257989
R7154 VB_A.n43 VB_A.n42 0.257989
R7155 VB_A.n44 VB_A.n43 0.257989
R7156 VB_A.n45 VB_A.n44 0.257989
R7157 VB_A.n46 VB_A.n45 0.257989
R7158 VB_A.n47 VB_A.n46 0.257989
R7159 VB_A.n48 VB_A.n47 0.257989
R7160 VB_A.n17 VB_A.n16 0.257989
R7161 VB_A.n18 VB_A.n17 0.257989
R7162 VB_A.n19 VB_A.n18 0.257989
R7163 VB_A.n20 VB_A.n19 0.257989
R7164 VB_A.n21 VB_A.n20 0.257989
R7165 VB_A.n22 VB_A.n21 0.257989
R7166 VB_A.n23 VB_A.n22 0.257989
R7167 VB_A.n24 VB_A.n23 0.257989
R7168 VB_A.n25 VB_A.n24 0.257989
R7169 VB_A.n26 VB_A.n25 0.257989
R7170 VB_A.n27 VB_A.n26 0.257989
R7171 VB_A.n28 VB_A.n27 0.257989
R7172 VB_A.n29 VB_A.n28 0.257989
R7173 VB_A.n30 VB_A.n29 0.257989
R7174 VB_A.n31 VB_A.n30 0.257989
R7175 VB_A.n1 VB_A.n0 0.257989
R7176 VB_A.n2 VB_A.n1 0.257989
R7177 VB_A.n3 VB_A.n2 0.257989
R7178 VB_A.n4 VB_A.n3 0.257989
R7179 VB_A.n5 VB_A.n4 0.257989
R7180 VB_A.n6 VB_A.n5 0.257989
R7181 VB_A.n7 VB_A.n6 0.257989
R7182 VB_A.n8 VB_A.n7 0.257989
R7183 VB_A.n9 VB_A.n8 0.257989
R7184 VB_A.n10 VB_A.n9 0.257989
R7185 VB_A.n11 VB_A.n10 0.257989
R7186 VB_A.n12 VB_A.n11 0.257989
R7187 VB_A.n13 VB_A.n12 0.257989
R7188 VB_A.n14 VB_A.n13 0.257989
R7189 VB_A.n15 VB_A.n14 0.257989
R7190 VB_A.n100 VB_A.n99 0.192994
R7191 VB_A.n83 VB_A.n82 0.192161
R7192 VB_A.n66 VB_A.n65 0.192161
R7193 VB_A.n49 VB_A.n48 0.192161
R7194 VB_A.n32 VB_A.n31 0.192161
R7195 IB.n22 IB.t12 22.9549
R7196 IB.n17 IB.t19 22.9549
R7197 IB.n12 IB.t22 22.9549
R7198 IB.n7 IB.t24 22.9549
R7199 IB.n27 IB.t33 22.9537
R7200 IB.n3 IB.t14 22.9537
R7201 IB.n27 IB.t20 22.5678
R7202 IB.n28 IB.t26 22.5678
R7203 IB.n29 IB.t32 22.5678
R7204 IB.n30 IB.t27 22.5678
R7205 IB.n22 IB.t17 22.5678
R7206 IB.n23 IB.t15 22.5678
R7207 IB.n24 IB.t31 22.5678
R7208 IB.n25 IB.t18 22.5678
R7209 IB.n17 IB.t4 22.5678
R7210 IB.n18 IB.t6 22.5678
R7211 IB.n19 IB.t8 22.5678
R7212 IB.n20 IB.t23 22.5678
R7213 IB.n12 IB.t0 22.5678
R7214 IB.n13 IB.t2 22.5678
R7215 IB.n14 IB.t11 22.5678
R7216 IB.n15 IB.t25 22.5678
R7217 IB.n7 IB.t30 22.5678
R7218 IB.n8 IB.t29 22.5678
R7219 IB.n9 IB.t16 22.5678
R7220 IB.n10 IB.t21 22.5678
R7221 IB.n3 IB.t28 22.5678
R7222 IB.n4 IB.t9 22.5678
R7223 IB.n5 IB.t13 22.5678
R7224 IB.n6 IB.t10 22.5678
R7225 IB.n0 IB.t3 5.71641
R7226 IB.n0 IB.t7 5.71641
R7227 IB.n1 IB.t1 5.71419
R7228 IB.n1 IB.t5 5.71419
R7229 IB.n32 IB.n2 2.42598
R7230 IB IB.n32 2.1409
R7231 IB.n2 IB.n1 0.844754
R7232 IB.n32 IB.n31 0.813
R7233 IB.n11 IB.n6 0.517817
R7234 IB.n10 IB.n9 0.390134
R7235 IB.n19 IB.n18 0.388884
R7236 IB.n14 IB.n13 0.388884
R7237 IB.n25 IB.n24 0.387009
R7238 IB.n28 IB.n27 0.386384
R7239 IB.n29 IB.n28 0.386384
R7240 IB.n30 IB.n29 0.386384
R7241 IB.n23 IB.n22 0.386384
R7242 IB.n24 IB.n23 0.386384
R7243 IB.n18 IB.n17 0.386384
R7244 IB.n20 IB.n19 0.386384
R7245 IB.n13 IB.n12 0.386384
R7246 IB.n15 IB.n14 0.386384
R7247 IB.n8 IB.n7 0.386384
R7248 IB.n9 IB.n8 0.386384
R7249 IB.n4 IB.n3 0.386384
R7250 IB.n5 IB.n4 0.386384
R7251 IB.n6 IB.n5 0.386384
R7252 IB.n31 IB.n30 0.267817
R7253 IB.n26 IB.n25 0.265942
R7254 IB.n21 IB.n20 0.264067
R7255 IB.n16 IB.n15 0.264067
R7256 IB.n11 IB.n10 0.262817
R7257 IB.n16 IB.n11 0.2505
R7258 IB.n21 IB.n16 0.2505
R7259 IB.n26 IB.n21 0.2505
R7260 IB.n31 IB.n26 0.2505
R7261 IB.n2 IB.n0 0.00820634
R7262 dummy_100.n8 dummy_100.t5 8.28993
R7263 dummy_100.n3 dummy_100.t32 8.13564
R7264 dummy_100.n2 dummy_100.t39 8.13411
R7265 dummy_100.n2 dummy_100.t24 5.71419
R7266 dummy_100.n2 dummy_100.t15 5.71419
R7267 dummy_100.n1 dummy_100.t25 5.71419
R7268 dummy_100.n1 dummy_100.t6 5.71419
R7269 dummy_100.n28 dummy_100.t2 5.71419
R7270 dummy_100.n29 dummy_100.t8 5.71419
R7271 dummy_100.n30 dummy_100.t20 5.71419
R7272 dummy_100.n31 dummy_100.t0 5.71419
R7273 dummy_100.n31 dummy_100.t31 5.71419
R7274 dummy_100.n15 dummy_100.t26 5.71419
R7275 dummy_100.n14 dummy_100.t4 5.71419
R7276 dummy_100.n13 dummy_100.t36 5.71419
R7277 dummy_100.n12 dummy_100.t28 5.71419
R7278 dummy_100.n11 dummy_100.t34 5.71419
R7279 dummy_100.n5 dummy_100.t11 5.71419
R7280 dummy_100.n5 dummy_100.t14 5.71419
R7281 dummy_100.n4 dummy_100.t33 5.71419
R7282 dummy_100.n4 dummy_100.t38 5.71419
R7283 dummy_100.n3 dummy_100.t10 5.71419
R7284 dummy_100.n3 dummy_100.t19 5.71419
R7285 dummy_100.n0 dummy_100.t35 5.71419
R7286 dummy_100.n0 dummy_100.t18 5.71419
R7287 dummy_100.n9 dummy_100.t29 5.71419
R7288 dummy_100.n8 dummy_100.t37 5.71419
R7289 dummy_100.n17 dummy_100.t12 5.71419
R7290 dummy_100.n17 dummy_100.t27 5.71419
R7291 dummy_100.n18 dummy_100.t16 5.71419
R7292 dummy_100.n18 dummy_100.t13 5.71419
R7293 dummy_100.n19 dummy_100.t22 5.71419
R7294 dummy_100.n19 dummy_100.t17 5.71419
R7295 dummy_100.n20 dummy_100.t30 5.71419
R7296 dummy_100.n20 dummy_100.t23 5.71419
R7297 dummy_100.n25 dummy_100.t1 5.71419
R7298 dummy_100.n24 dummy_100.t21 5.71419
R7299 dummy_100.n23 dummy_100.t9 5.71419
R7300 dummy_100.n22 dummy_100.t3 5.71419
R7301 dummy_100.n21 dummy_100.t7 5.71419
R7302 dummy_100.n11 dummy_100.n10 5.02967
R7303 dummy_100.n32 dummy_100.n25 3.91962
R7304 dummy_100.n12 dummy_100.n11 2.82133
R7305 dummy_100.n13 dummy_100.n12 2.82133
R7306 dummy_100.n14 dummy_100.n13 2.82133
R7307 dummy_100.n15 dummy_100.n14 2.82133
R7308 dummy_100.n30 dummy_100.n29 2.82133
R7309 dummy_100.n29 dummy_100.n28 2.82133
R7310 dummy_100.n9 dummy_100.n8 2.57624
R7311 dummy_100.n22 dummy_100.n21 2.57624
R7312 dummy_100.n23 dummy_100.n22 2.57624
R7313 dummy_100.n24 dummy_100.n23 2.57624
R7314 dummy_100.n25 dummy_100.n24 2.57624
R7315 dummy_100.n28 dummy_100.n1 2.13481
R7316 dummy_100.n31 dummy_100.n30 2.11211
R7317 dummy_100.n7 dummy_100.n6 2.063
R7318 dummy_100.n10 dummy_100.n7 2.063
R7319 dummy_100 dummy_100.n36 2.063
R7320 dummy_100.n36 dummy_100.n35 2.063
R7321 dummy_100.n35 dummy_100.n34 2.063
R7322 dummy_100.n34 dummy_100.n33 2.063
R7323 dummy_100.n33 dummy_100.n32 2.063
R7324 dummy_100.n27 dummy_100.n26 2.063
R7325 dummy_100.n0 dummy_100.n9 2.00834
R7326 dummy_100.n16 dummy_100.n15 1.91717
R7327 dummy_100.n7 dummy_100.n3 1.30616
R7328 dummy_100.n26 dummy_100.n2 1.1639
R7329 dummy_100.n1 dummy_100.n27 1.08801
R7330 dummy_100.n10 dummy_100.n0 0.881161
R7331 dummy_100.n5 dummy_100.n4 0.876108
R7332 dummy_100.n6 dummy_100.n5 0.872233
R7333 dummy_100.n36 dummy_100.n17 0.600804
R7334 dummy_100.n35 dummy_100.n18 0.600804
R7335 dummy_100.n34 dummy_100.n19 0.600804
R7336 dummy_100.n33 dummy_100.n20 0.600804
R7337 dummy_100.n32 dummy_100.n31 0.600804
R7338 dummy_100.n16 dummy_100 0.1255
R7339 dummy_100 dummy_100.n16 0.063
R7340 dummy_3.n28 dummy_3.t19 4.44742
R7341 dummy_3.n60 dummy_3.t20 4.42883
R7342 dummy_3.n2 dummy_3.t14 3.52072
R7343 dummy_3.n11 dummy_3.t13 3.51909
R7344 dummy_3.n4 dummy_3.t6 3.51864
R7345 dummy_3.n6 dummy_3.t82 3.51864
R7346 dummy_3.n8 dummy_3.t74 3.51864
R7347 dummy_3.n10 dummy_3.t16 3.51864
R7348 dummy_3.n7 dummy_3.t75 3.51707
R7349 dummy_3.n3 dummy_3.t7 3.51707
R7350 dummy_3.n9 dummy_3.t17 3.51707
R7351 dummy_3.n5 dummy_3.t83 3.51558
R7352 dummy_3.n83 dummy_3.t50 3.48747
R7353 dummy_3.n81 dummy_3.t10 3.48747
R7354 dummy_3.n79 dummy_3.t62 3.48747
R7355 dummy_3.n77 dummy_3.t22 3.48747
R7356 dummy_3.n82 dummy_3.t51 3.4869
R7357 dummy_3.n78 dummy_3.t63 3.4869
R7358 dummy_3.n76 dummy_3.t23 3.4869
R7359 dummy_3.n80 dummy_3.t11 3.48662
R7360 dummy_3.n84 dummy_3.t38 3.48393
R7361 dummy_3.n74 dummy_3.t76 3.48239
R7362 dummy_3.n1 dummy_3.t15 3.48239
R7363 dummy_3.n12 dummy_3.t12 3.48239
R7364 dummy_3.n59 dummy_3.t77 3.48239
R7365 dummy_3.n44 dummy_3.t21 3.48118
R7366 dummy_3.n45 dummy_3.t47 3.48118
R7367 dummy_3.n46 dummy_3.t61 3.48118
R7368 dummy_3.n47 dummy_3.t71 3.48118
R7369 dummy_3.n48 dummy_3.t41 3.48118
R7370 dummy_3.n49 dummy_3.t53 3.48118
R7371 dummy_3.n50 dummy_3.t27 3.48118
R7372 dummy_3.n51 dummy_3.t31 3.48118
R7373 dummy_3.n52 dummy_3.t35 3.48118
R7374 dummy_3.n53 dummy_3.t3 3.48118
R7375 dummy_3.n54 dummy_3.t9 3.48118
R7376 dummy_3.n55 dummy_3.t79 3.48118
R7377 dummy_3.n56 dummy_3.t81 3.48118
R7378 dummy_3.n57 dummy_3.t1 3.48118
R7379 dummy_3.n58 dummy_3.t5 3.48118
R7380 dummy_3.n73 dummy_3.t4 3.48118
R7381 dummy_3.n72 dummy_3.t0 3.48118
R7382 dummy_3.n71 dummy_3.t80 3.48118
R7383 dummy_3.n70 dummy_3.t78 3.48118
R7384 dummy_3.n69 dummy_3.t8 3.48118
R7385 dummy_3.n68 dummy_3.t2 3.48118
R7386 dummy_3.n67 dummy_3.t34 3.48118
R7387 dummy_3.n66 dummy_3.t30 3.48118
R7388 dummy_3.n65 dummy_3.t26 3.48118
R7389 dummy_3.n64 dummy_3.t52 3.48118
R7390 dummy_3.n63 dummy_3.t40 3.48118
R7391 dummy_3.n62 dummy_3.t70 3.48118
R7392 dummy_3.n61 dummy_3.t60 3.48118
R7393 dummy_3.n60 dummy_3.t46 3.48118
R7394 dummy_3.n41 dummy_3.t69 3.48118
R7395 dummy_3.n40 dummy_3.t59 3.48118
R7396 dummy_3.n39 dummy_3.t55 3.48118
R7397 dummy_3.n38 dummy_3.t45 3.48118
R7398 dummy_3.n37 dummy_3.t73 3.48118
R7399 dummy_3.n36 dummy_3.t65 3.48118
R7400 dummy_3.n35 dummy_3.t33 3.48118
R7401 dummy_3.n34 dummy_3.t29 3.48118
R7402 dummy_3.n33 dummy_3.t25 3.48118
R7403 dummy_3.n32 dummy_3.t49 3.48118
R7404 dummy_3.n31 dummy_3.t37 3.48118
R7405 dummy_3.n30 dummy_3.t67 3.48118
R7406 dummy_3.n29 dummy_3.t57 3.48118
R7407 dummy_3.n28 dummy_3.t43 3.48118
R7408 dummy_3.n27 dummy_3.t68 3.48118
R7409 dummy_3.n26 dummy_3.t58 3.48118
R7410 dummy_3.n25 dummy_3.t54 3.48118
R7411 dummy_3.n24 dummy_3.t44 3.48118
R7412 dummy_3.n23 dummy_3.t72 3.48118
R7413 dummy_3.n22 dummy_3.t64 3.48118
R7414 dummy_3.n21 dummy_3.t32 3.48118
R7415 dummy_3.n20 dummy_3.t28 3.48118
R7416 dummy_3.n19 dummy_3.t24 3.48118
R7417 dummy_3.n18 dummy_3.t48 3.48118
R7418 dummy_3.n17 dummy_3.t36 3.48118
R7419 dummy_3.n16 dummy_3.t66 3.48118
R7420 dummy_3.n15 dummy_3.t56 3.48118
R7421 dummy_3.n14 dummy_3.t42 3.48118
R7422 dummy_3.n13 dummy_3.t18 3.48118
R7423 dummy_3.n0 dummy_3.t39 3.48093
R7424 dummy_3.n43 dummy_3.n41 1.44478
R7425 dummy_3.n29 dummy_3.n28 0.966748
R7426 dummy_3.n30 dummy_3.n29 0.966748
R7427 dummy_3.n31 dummy_3.n30 0.966748
R7428 dummy_3.n32 dummy_3.n31 0.966748
R7429 dummy_3.n33 dummy_3.n32 0.966748
R7430 dummy_3.n34 dummy_3.n33 0.966748
R7431 dummy_3.n35 dummy_3.n34 0.966748
R7432 dummy_3.n36 dummy_3.n35 0.966748
R7433 dummy_3.n37 dummy_3.n36 0.966748
R7434 dummy_3.n38 dummy_3.n37 0.966748
R7435 dummy_3.n39 dummy_3.n38 0.966748
R7436 dummy_3.n40 dummy_3.n39 0.966748
R7437 dummy_3.n41 dummy_3.n40 0.966748
R7438 dummy_3.n58 dummy_3.n57 0.966748
R7439 dummy_3.n57 dummy_3.n56 0.966748
R7440 dummy_3.n56 dummy_3.n55 0.966748
R7441 dummy_3.n55 dummy_3.n54 0.966748
R7442 dummy_3.n54 dummy_3.n53 0.966748
R7443 dummy_3.n53 dummy_3.n52 0.966748
R7444 dummy_3.n52 dummy_3.n51 0.966748
R7445 dummy_3.n51 dummy_3.n50 0.966748
R7446 dummy_3.n50 dummy_3.n49 0.966748
R7447 dummy_3.n49 dummy_3.n48 0.966748
R7448 dummy_3.n48 dummy_3.n47 0.966748
R7449 dummy_3.n47 dummy_3.n46 0.966748
R7450 dummy_3.n46 dummy_3.n45 0.966748
R7451 dummy_3.n45 dummy_3.n44 0.966748
R7452 dummy_3.n61 dummy_3.n60 0.948155
R7453 dummy_3.n62 dummy_3.n61 0.948155
R7454 dummy_3.n63 dummy_3.n62 0.948155
R7455 dummy_3.n64 dummy_3.n63 0.948155
R7456 dummy_3.n65 dummy_3.n64 0.948155
R7457 dummy_3.n66 dummy_3.n65 0.948155
R7458 dummy_3.n67 dummy_3.n66 0.948155
R7459 dummy_3.n68 dummy_3.n67 0.948155
R7460 dummy_3.n69 dummy_3.n68 0.948155
R7461 dummy_3.n70 dummy_3.n69 0.948155
R7462 dummy_3.n71 dummy_3.n70 0.948155
R7463 dummy_3.n72 dummy_3.n71 0.948155
R7464 dummy_3.n73 dummy_3.n72 0.948155
R7465 dummy_3.n14 dummy_3.n13 0.948155
R7466 dummy_3.n15 dummy_3.n14 0.948155
R7467 dummy_3.n16 dummy_3.n15 0.948155
R7468 dummy_3.n17 dummy_3.n16 0.948155
R7469 dummy_3.n18 dummy_3.n17 0.948155
R7470 dummy_3.n19 dummy_3.n18 0.948155
R7471 dummy_3.n20 dummy_3.n19 0.948155
R7472 dummy_3.n21 dummy_3.n20 0.948155
R7473 dummy_3.n22 dummy_3.n21 0.948155
R7474 dummy_3.n23 dummy_3.n22 0.948155
R7475 dummy_3.n24 dummy_3.n23 0.948155
R7476 dummy_3.n25 dummy_3.n24 0.948155
R7477 dummy_3.n26 dummy_3.n25 0.948155
R7478 dummy_3.n27 dummy_3.n26 0.948155
R7479 dummy_3.n59 dummy_3.n58 0.909211
R7480 dummy_3.n13 dummy_3.n12 0.898657
R7481 dummy_3.n74 dummy_3.n73 0.894942
R7482 dummy_3 dummy_3.n27 0.489506
R7483 dummy_3 dummy_3.n84 0.40075
R7484 dummy_3.n12 dummy_3.n11 0.334804
R7485 dummy_3.n2 dummy_3.n1 0.334348
R7486 dummy_3.n75 dummy_3.n59 0.326028
R7487 dummy_3.n6 dummy_3.n5 0.315662
R7488 dummy_3.n83 dummy_3.n82 0.315161
R7489 dummy_3.n79 dummy_3.n78 0.315161
R7490 dummy_3.n77 dummy_3.n76 0.315161
R7491 dummy_3.n10 dummy_3.n9 0.315161
R7492 dummy_3.n4 dummy_3.n3 0.315161
R7493 dummy_3.n8 dummy_3.n7 0.315161
R7494 dummy_3.n84 dummy_3.n0 0.314676
R7495 dummy_3.n81 dummy_3.n80 0.311871
R7496 dummy_3.n80 dummy_3.n79 0.150815
R7497 dummy_3.n7 dummy_3.n6 0.147546
R7498 dummy_3.n3 dummy_3.n2 0.141668
R7499 dummy_3.n76 dummy_3.n75 0.141275
R7500 dummy_3.n82 dummy_3.n81 0.141045
R7501 dummy_3.n78 dummy_3.n77 0.141045
R7502 dummy_3.n11 dummy_3.n10 0.141045
R7503 dummy_3.n9 dummy_3.n8 0.141045
R7504 dummy_3.n5 dummy_3.n4 0.140588
R7505 dummy_3.n0 dummy_3.n83 0.104757
R7506 dummy_3.n0 dummy_3.n43 0.0932417
R7507 dummy_3.n43 dummy_3.n42 0.0377984
R7508 dummy_3.n75 dummy_3.n74 0.0118634
R7509 dummy_2.n21 dummy_2.t2 5.78964
R7510 dummy_2.n20 dummy_2.t3 5.7861
R7511 dummy_2.n23 dummy_2.t36 5.7826
R7512 dummy_2.n25 dummy_2.t70 5.77927
R7513 dummy_2.n24 dummy_2.t71 5.77101
R7514 dummy_2.n27 dummy_2.t26 5.76803
R7515 dummy_2.n26 dummy_2.t27 5.76437
R7516 dummy_2.n22 dummy_2.t37 5.76437
R7517 dummy_2.n61 dummy_2.t33 5.72689
R7518 dummy_2.n83 dummy_2.t11 5.72634
R7519 dummy_2.n82 dummy_2.t54 5.72583
R7520 dummy_2.n84 dummy_2.t10 5.72583
R7521 dummy_2.n80 dummy_2.t20 5.7255
R7522 dummy_2.n79 dummy_2.t21 5.72533
R7523 dummy_2.n81 dummy_2.t55 5.72533
R7524 dummy_2.n78 dummy_2.t72 5.72477
R7525 dummy_2.n77 dummy_2.t73 5.72455
R7526 dummy_2.n0 dummy_2.t9 5.72347
R7527 dummy_2.n85 dummy_2.t8 5.72347
R7528 dummy_2.n1 dummy_2.t32 5.72247
R7529 dummy_2.n29 dummy_2.t79 5.7154
R7530 dummy_2.n45 dummy_2.t17 5.7154
R7531 dummy_2.n2 dummy_2.t78 5.7154
R7532 dummy_2.n18 dummy_2.t16 5.7154
R7533 dummy_2.n49 dummy_2.t39 5.71419
R7534 dummy_2.n50 dummy_2.t81 5.71419
R7535 dummy_2.n51 dummy_2.t1 5.71419
R7536 dummy_2.n52 dummy_2.t67 5.71419
R7537 dummy_2.n53 dummy_2.t25 5.71419
R7538 dummy_2.n54 dummy_2.t65 5.71419
R7539 dummy_2.n55 dummy_2.t51 5.71419
R7540 dummy_2.n56 dummy_2.t69 5.71419
R7541 dummy_2.n57 dummy_2.t49 5.71419
R7542 dummy_2.n58 dummy_2.t31 5.71419
R7543 dummy_2.n59 dummy_2.t13 5.71419
R7544 dummy_2.n60 dummy_2.t77 5.71419
R7545 dummy_2.n76 dummy_2.t76 5.71419
R7546 dummy_2.n75 dummy_2.t12 5.71419
R7547 dummy_2.n74 dummy_2.t30 5.71419
R7548 dummy_2.n73 dummy_2.t48 5.71419
R7549 dummy_2.n72 dummy_2.t68 5.71419
R7550 dummy_2.n71 dummy_2.t50 5.71419
R7551 dummy_2.n70 dummy_2.t64 5.71419
R7552 dummy_2.n69 dummy_2.t24 5.71419
R7553 dummy_2.n68 dummy_2.t66 5.71419
R7554 dummy_2.n67 dummy_2.t0 5.71419
R7555 dummy_2.n66 dummy_2.t80 5.71419
R7556 dummy_2.n65 dummy_2.t38 5.71419
R7557 dummy_2.n64 dummy_2.t82 5.71419
R7558 dummy_2.n63 dummy_2.t40 5.71419
R7559 dummy_2.n62 dummy_2.t56 5.71419
R7560 dummy_2.n3 dummy_2.t34 5.71419
R7561 dummy_2.n4 dummy_2.t18 5.71419
R7562 dummy_2.n5 dummy_2.t60 5.71419
R7563 dummy_2.n6 dummy_2.t14 5.71419
R7564 dummy_2.n7 dummy_2.t58 5.71419
R7565 dummy_2.n8 dummy_2.t62 5.71419
R7566 dummy_2.n9 dummy_2.t44 5.71419
R7567 dummy_2.n10 dummy_2.t4 5.71419
R7568 dummy_2.n11 dummy_2.t42 5.71419
R7569 dummy_2.n12 dummy_2.t28 5.71419
R7570 dummy_2.n13 dummy_2.t46 5.71419
R7571 dummy_2.n14 dummy_2.t22 5.71419
R7572 dummy_2.n15 dummy_2.t6 5.71419
R7573 dummy_2.n16 dummy_2.t74 5.71419
R7574 dummy_2.n17 dummy_2.t52 5.71419
R7575 dummy_2.n30 dummy_2.t35 5.71419
R7576 dummy_2.n31 dummy_2.t19 5.71419
R7577 dummy_2.n32 dummy_2.t61 5.71419
R7578 dummy_2.n33 dummy_2.t15 5.71419
R7579 dummy_2.n34 dummy_2.t59 5.71419
R7580 dummy_2.n35 dummy_2.t63 5.71419
R7581 dummy_2.n36 dummy_2.t45 5.71419
R7582 dummy_2.n37 dummy_2.t5 5.71419
R7583 dummy_2.n38 dummy_2.t43 5.71419
R7584 dummy_2.n39 dummy_2.t29 5.71419
R7585 dummy_2.n40 dummy_2.t47 5.71419
R7586 dummy_2.n41 dummy_2.t23 5.71419
R7587 dummy_2.n42 dummy_2.t7 5.71419
R7588 dummy_2.n43 dummy_2.t75 5.71419
R7589 dummy_2.n44 dummy_2.t53 5.71419
R7590 dummy_2.n46 dummy_2.t57 5.71419
R7591 dummy_2.n47 dummy_2.t41 5.71419
R7592 dummy_2.n48 dummy_2.t83 5.71419
R7593 dummy_2.n17 dummy_2.n16 1.61925
R7594 dummy_2.n16 dummy_2.n15 1.61925
R7595 dummy_2.n15 dummy_2.n14 1.61925
R7596 dummy_2.n14 dummy_2.n13 1.61925
R7597 dummy_2.n13 dummy_2.n12 1.61925
R7598 dummy_2.n12 dummy_2.n11 1.61925
R7599 dummy_2.n11 dummy_2.n10 1.61925
R7600 dummy_2.n10 dummy_2.n9 1.61925
R7601 dummy_2.n9 dummy_2.n8 1.61925
R7602 dummy_2.n8 dummy_2.n7 1.61925
R7603 dummy_2.n7 dummy_2.n6 1.61925
R7604 dummy_2.n6 dummy_2.n5 1.61925
R7605 dummy_2.n5 dummy_2.n4 1.61925
R7606 dummy_2.n4 dummy_2.n3 1.61925
R7607 dummy_2.n63 dummy_2.n62 1.61925
R7608 dummy_2.n64 dummy_2.n63 1.61925
R7609 dummy_2.n65 dummy_2.n64 1.61925
R7610 dummy_2.n66 dummy_2.n65 1.61925
R7611 dummy_2.n67 dummy_2.n66 1.61925
R7612 dummy_2.n68 dummy_2.n67 1.61925
R7613 dummy_2.n69 dummy_2.n68 1.61925
R7614 dummy_2.n70 dummy_2.n69 1.61925
R7615 dummy_2.n71 dummy_2.n70 1.61925
R7616 dummy_2.n72 dummy_2.n71 1.61925
R7617 dummy_2.n73 dummy_2.n72 1.61925
R7618 dummy_2.n74 dummy_2.n73 1.61925
R7619 dummy_2.n75 dummy_2.n74 1.61925
R7620 dummy_2.n76 dummy_2.n75 1.61925
R7621 dummy_2.n3 dummy_2.n2 1.5435
R7622 dummy_2.n44 dummy_2.n43 1.52666
R7623 dummy_2.n43 dummy_2.n42 1.52666
R7624 dummy_2.n42 dummy_2.n41 1.52666
R7625 dummy_2.n41 dummy_2.n40 1.52666
R7626 dummy_2.n40 dummy_2.n39 1.52666
R7627 dummy_2.n39 dummy_2.n38 1.52666
R7628 dummy_2.n38 dummy_2.n37 1.52666
R7629 dummy_2.n37 dummy_2.n36 1.52666
R7630 dummy_2.n36 dummy_2.n35 1.52666
R7631 dummy_2.n35 dummy_2.n34 1.52666
R7632 dummy_2.n34 dummy_2.n33 1.52666
R7633 dummy_2.n33 dummy_2.n32 1.52666
R7634 dummy_2.n32 dummy_2.n31 1.52666
R7635 dummy_2.n31 dummy_2.n30 1.52666
R7636 dummy_2.n48 dummy_2.n47 1.52666
R7637 dummy_2.n47 dummy_2.n46 1.52666
R7638 dummy_2.n60 dummy_2.n59 1.52666
R7639 dummy_2.n59 dummy_2.n58 1.52666
R7640 dummy_2.n58 dummy_2.n57 1.52666
R7641 dummy_2.n57 dummy_2.n56 1.52666
R7642 dummy_2.n56 dummy_2.n55 1.52666
R7643 dummy_2.n55 dummy_2.n54 1.52666
R7644 dummy_2.n54 dummy_2.n53 1.52666
R7645 dummy_2.n53 dummy_2.n52 1.52666
R7646 dummy_2.n52 dummy_2.n51 1.52666
R7647 dummy_2.n51 dummy_2.n50 1.52666
R7648 dummy_2.n50 dummy_2.n49 1.52666
R7649 dummy_2.n49 dummy_2.n48 1.52666
R7650 dummy_2.n1 dummy_2.n76 1.49501
R7651 dummy_2.n30 dummy_2.n29 1.45576
R7652 dummy_2.n46 dummy_2.n45 1.45074
R7653 dummy_2.n0 dummy_2.n44 1.42
R7654 dummy_2.n61 dummy_2.n60 1.37201
R7655 dummy_2 dummy_2.n17 0.9005
R7656 dummy_2 dummy_2.n85 0.594012
R7657 dummy_2.n21 dummy_2.n20 0.315613
R7658 dummy_2.n85 dummy_2.n0 0.311881
R7659 dummy_2.n84 dummy_2.n83 0.309043
R7660 dummy_2.n82 dummy_2.n81 0.305753
R7661 dummy_2.n1 dummy_2.n61 0.30301
R7662 dummy_2.n25 dummy_2.n24 0.302464
R7663 dummy_2.n23 dummy_2.n22 0.302003
R7664 dummy_2.n80 dummy_2.n79 0.298714
R7665 dummy_2.n27 dummy_2.n26 0.295424
R7666 dummy_2.n78 dummy_2.n77 0.292135
R7667 dummy_2.n79 dummy_2.n78 0.163912
R7668 dummy_2.n28 dummy_2.n27 0.160656
R7669 dummy_2.n81 dummy_2.n80 0.160656
R7670 dummy_2.n77 dummy_2.n1 0.158896
R7671 dummy_2.n24 dummy_2.n23 0.157389
R7672 dummy_2.n20 dummy_2.n19 0.154555
R7673 dummy_2.n26 dummy_2.n25 0.140127
R7674 dummy_2.n22 dummy_2.n21 0.140114
R7675 dummy_2.n83 dummy_2.n82 0.133605
R7676 dummy_2.n0 dummy_2.n84 0.131394
R7677 dummy_2.n19 dummy_2.n18 0.0421669
R7678 dummy_2.n29 dummy_2.n28 0.0421635
R7679 OUT.n42 OUT.t0 6.70615
R7680 OUT.n14 OUT.t21 6.66895
R7681 OUT.n56 OUT.n55 6.62597
R7682 OUT.n57 OUT.n27 6.44828
R7683 OUT.n55 OUT.t2 5.71419
R7684 OUT.n54 OUT.t25 5.71419
R7685 OUT.n53 OUT.t3 5.71419
R7686 OUT.n52 OUT.t24 5.71419
R7687 OUT.n51 OUT.t11 5.71419
R7688 OUT.n50 OUT.t14 5.71419
R7689 OUT.n49 OUT.t8 5.71419
R7690 OUT.n48 OUT.t12 5.71419
R7691 OUT.n47 OUT.t7 5.71419
R7692 OUT.n46 OUT.t19 5.71419
R7693 OUT.n45 OUT.t9 5.71419
R7694 OUT.n44 OUT.t29 5.71419
R7695 OUT.n43 OUT.t15 5.71419
R7696 OUT.n42 OUT.t16 5.71419
R7697 OUT.n27 OUT.t22 5.71419
R7698 OUT.n26 OUT.t18 5.71419
R7699 OUT.n25 OUT.t23 5.71419
R7700 OUT.n24 OUT.t17 5.71419
R7701 OUT.n23 OUT.t1 5.71419
R7702 OUT.n22 OUT.t5 5.71419
R7703 OUT.n21 OUT.t27 5.71419
R7704 OUT.n20 OUT.t4 5.71419
R7705 OUT.n19 OUT.t26 5.71419
R7706 OUT.n18 OUT.t13 5.71419
R7707 OUT.n17 OUT.t28 5.71419
R7708 OUT.n16 OUT.t20 5.71419
R7709 OUT.n15 OUT.t6 5.71419
R7710 OUT.n14 OUT.t10 5.71419
R7711 OUT.n56 OUT.n41 5.60595
R7712 OUT.n28 OUT.t42 4.44742
R7713 OUT.n0 OUT.t54 4.42883
R7714 OUT.n58 OUT.n13 3.96778
R7715 OUT.n13 OUT.t59 3.48118
R7716 OUT.n12 OUT.t56 3.48118
R7717 OUT.n11 OUT.t52 3.48118
R7718 OUT.n10 OUT.t31 3.48118
R7719 OUT.n9 OUT.t41 3.48118
R7720 OUT.n8 OUT.t55 3.48118
R7721 OUT.n7 OUT.t43 3.48118
R7722 OUT.n6 OUT.t50 3.48118
R7723 OUT.n5 OUT.t47 3.48118
R7724 OUT.n4 OUT.t35 3.48118
R7725 OUT.n3 OUT.t53 3.48118
R7726 OUT.n2 OUT.t30 3.48118
R7727 OUT.n1 OUT.t32 3.48118
R7728 OUT.n0 OUT.t36 3.48118
R7729 OUT.n41 OUT.t34 3.48118
R7730 OUT.n40 OUT.t45 3.48118
R7731 OUT.n39 OUT.t37 3.48118
R7732 OUT.n38 OUT.t38 3.48118
R7733 OUT.n37 OUT.t48 3.48118
R7734 OUT.n36 OUT.t46 3.48118
R7735 OUT.n35 OUT.t51 3.48118
R7736 OUT.n34 OUT.t44 3.48118
R7737 OUT.n33 OUT.t57 3.48118
R7738 OUT.n32 OUT.t33 3.48118
R7739 OUT.n31 OUT.t49 3.48118
R7740 OUT.n30 OUT.t58 3.48118
R7741 OUT.n29 OUT.t39 3.48118
R7742 OUT.n28 OUT.t40 3.48118
R7743 OUT OUT.n58 2.8909
R7744 OUT.n57 OUT.n56 1.53459
R7745 OUT.n43 OUT.n42 0.992464
R7746 OUT.n44 OUT.n43 0.992464
R7747 OUT.n45 OUT.n44 0.992464
R7748 OUT.n46 OUT.n45 0.992464
R7749 OUT.n47 OUT.n46 0.992464
R7750 OUT.n48 OUT.n47 0.992464
R7751 OUT.n49 OUT.n48 0.992464
R7752 OUT.n50 OUT.n49 0.992464
R7753 OUT.n51 OUT.n50 0.992464
R7754 OUT.n52 OUT.n51 0.992464
R7755 OUT.n53 OUT.n52 0.992464
R7756 OUT.n54 OUT.n53 0.992464
R7757 OUT.n55 OUT.n54 0.992464
R7758 OUT.n29 OUT.n28 0.966748
R7759 OUT.n30 OUT.n29 0.966748
R7760 OUT.n31 OUT.n30 0.966748
R7761 OUT.n32 OUT.n31 0.966748
R7762 OUT.n33 OUT.n32 0.966748
R7763 OUT.n34 OUT.n33 0.966748
R7764 OUT.n35 OUT.n34 0.966748
R7765 OUT.n36 OUT.n35 0.966748
R7766 OUT.n37 OUT.n36 0.966748
R7767 OUT.n38 OUT.n37 0.966748
R7768 OUT.n39 OUT.n38 0.966748
R7769 OUT.n40 OUT.n39 0.966748
R7770 OUT.n41 OUT.n40 0.966748
R7771 OUT.n15 OUT.n14 0.955262
R7772 OUT.n16 OUT.n15 0.955262
R7773 OUT.n17 OUT.n16 0.955262
R7774 OUT.n18 OUT.n17 0.955262
R7775 OUT.n19 OUT.n18 0.955262
R7776 OUT.n20 OUT.n19 0.955262
R7777 OUT.n21 OUT.n20 0.955262
R7778 OUT.n22 OUT.n21 0.955262
R7779 OUT.n23 OUT.n22 0.955262
R7780 OUT.n24 OUT.n23 0.955262
R7781 OUT.n25 OUT.n24 0.955262
R7782 OUT.n26 OUT.n25 0.955262
R7783 OUT.n27 OUT.n26 0.955262
R7784 OUT.n1 OUT.n0 0.948155
R7785 OUT.n2 OUT.n1 0.948155
R7786 OUT.n3 OUT.n2 0.948155
R7787 OUT.n4 OUT.n3 0.948155
R7788 OUT.n5 OUT.n4 0.948155
R7789 OUT.n6 OUT.n5 0.948155
R7790 OUT.n7 OUT.n6 0.948155
R7791 OUT.n8 OUT.n7 0.948155
R7792 OUT.n9 OUT.n8 0.948155
R7793 OUT.n10 OUT.n9 0.948155
R7794 OUT.n11 OUT.n10 0.948155
R7795 OUT.n12 OUT.n11 0.948155
R7796 OUT.n13 OUT.n12 0.948155
R7797 OUT.n58 OUT.n57 0.606899
R7798 IN_M.n107 IN_M.t15 746.848
R7799 IN_M.n121 IN_M.t0 746.846
R7800 IN_M.n120 IN_M.t9 746.846
R7801 IN_M.n119 IN_M.t10 746.846
R7802 IN_M.n118 IN_M.t23 746.846
R7803 IN_M.n117 IN_M.t29 746.846
R7804 IN_M.n116 IN_M.t21 746.846
R7805 IN_M.n115 IN_M.t26 746.846
R7806 IN_M.n114 IN_M.t16 746.846
R7807 IN_M.n113 IN_M.t27 746.846
R7808 IN_M.n112 IN_M.t2 746.846
R7809 IN_M.n111 IN_M.t3 746.846
R7810 IN_M.n110 IN_M.t20 746.846
R7811 IN_M.n217 IN_M.t4 746.846
R7812 IN_M.n0 IN_M.t24 746.846
R7813 IN_M.n1 IN_M.t14 746.846
R7814 IN_M.n2 IN_M.t13 746.846
R7815 IN_M.n3 IN_M.t6 746.846
R7816 IN_M.n4 IN_M.t22 746.846
R7817 IN_M.n5 IN_M.t5 746.846
R7818 IN_M.n6 IN_M.t25 746.846
R7819 IN_M.n8 IN_M.t28 746.846
R7820 IN_M.n9 IN_M.t18 746.846
R7821 IN_M.n10 IN_M.t17 746.846
R7822 IN_M.n11 IN_M.t8 746.846
R7823 IN_M.n122 IN_M.t12 746.309
R7824 IN_M.n7 IN_M.t7 746.309
R7825 IN_M.n12 IN_M.t19 746.309
R7826 IN_M.n123 IN_M.t1 374.077
R7827 IN_M.n13 IN_M.t11 374.077
R7828 IN_M IN_M.n220 4.0484
R7829 IN_M.n220 IN_M.n219 3.00474
R7830 IN_M.n220 IN_M.n109 2.85474
R7831 IN_M.n124 IN_M.n123 2.43766
R7832 IN_M.n14 IN_M.n13 2.43766
R7833 IN_M.n49 IN_M.n48 2.35675
R7834 IN_M.n159 IN_M.n158 2.34135
R7835 IN_M.n166 IN_M.n165 2.33827
R7836 IN_M.n201 IN_M.n200 2.33827
R7837 IN_M.n91 IN_M.n90 2.33827
R7838 IN_M.n152 IN_M.n151 2.33055
R7839 IN_M.n145 IN_M.n144 2.32981
R7840 IN_M.n180 IN_M.n179 2.32981
R7841 IN_M.n35 IN_M.n34 2.32981
R7842 IN_M.n70 IN_M.n69 2.32981
R7843 IN_M.n138 IN_M.n137 2.32981
R7844 IN_M.n173 IN_M.n172 2.32981
R7845 IN_M.n208 IN_M.n207 2.32981
R7846 IN_M.n28 IN_M.n27 2.32981
R7847 IN_M.n63 IN_M.n62 2.32981
R7848 IN_M.n98 IN_M.n97 2.32981
R7849 IN_M.n187 IN_M.n186 2.3298
R7850 IN_M.n42 IN_M.n41 2.3298
R7851 IN_M.n77 IN_M.n76 2.3298
R7852 IN_M.n194 IN_M.n193 2.32516
R7853 IN_M.n84 IN_M.n83 2.32442
R7854 IN_M.n131 IN_M.n130 2.32441
R7855 IN_M.n21 IN_M.n20 2.32441
R7856 IN_M.n56 IN_M.n55 2.32441
R7857 IN_M.n215 IN_M.n214 2.31935
R7858 IN_M.n105 IN_M.n104 2.29822
R7859 IN_M.n144 IN_M.n143 0.1243
R7860 IN_M.n179 IN_M.n178 0.1243
R7861 IN_M.n214 IN_M.n213 0.1243
R7862 IN_M.n34 IN_M.n33 0.1243
R7863 IN_M.n69 IN_M.n68 0.1243
R7864 IN_M.n104 IN_M.n103 0.1243
R7865 IN_M.n146 IN_M.n145 0.123792
R7866 IN_M.n181 IN_M.n180 0.123792
R7867 IN_M.n36 IN_M.n35 0.123792
R7868 IN_M.n71 IN_M.n70 0.123792
R7869 IN_M.n137 IN_M.n136 0.123283
R7870 IN_M.n172 IN_M.n171 0.123283
R7871 IN_M.n207 IN_M.n206 0.123283
R7872 IN_M.n27 IN_M.n26 0.123283
R7873 IN_M.n62 IN_M.n61 0.123283
R7874 IN_M.n97 IN_M.n96 0.123283
R7875 IN_M.n188 IN_M.n187 0.122774
R7876 IN_M.n78 IN_M.n77 0.122774
R7877 IN_M.n151 IN_M.n150 0.121147
R7878 IN_M.n186 IN_M.n185 0.121147
R7879 IN_M.n41 IN_M.n40 0.121147
R7880 IN_M.n76 IN_M.n75 0.121147
R7881 IN_M.n139 IN_M.n138 0.120641
R7882 IN_M.n174 IN_M.n173 0.120641
R7883 IN_M.n209 IN_M.n208 0.120641
R7884 IN_M.n29 IN_M.n28 0.120641
R7885 IN_M.n64 IN_M.n63 0.120641
R7886 IN_M.n99 IN_M.n98 0.120641
R7887 IN_M.n153 IN_M.n152 0.114687
R7888 IN_M.n43 IN_M.n42 0.11444
R7889 IN_M.n193 IN_M.n192 0.113826
R7890 IN_M.n83 IN_M.n82 0.113826
R7891 IN_M.n132 IN_M.n131 0.11332
R7892 IN_M.n167 IN_M.n166 0.11332
R7893 IN_M.n202 IN_M.n201 0.11332
R7894 IN_M.n22 IN_M.n21 0.11332
R7895 IN_M.n57 IN_M.n56 0.11332
R7896 IN_M.n92 IN_M.n91 0.11332
R7897 IN_M.n165 IN_M.n164 0.113
R7898 IN_M.n200 IN_M.n199 0.113
R7899 IN_M.n90 IN_M.n89 0.113
R7900 IN_M.n125 IN_M.n124 0.110917
R7901 IN_M.n15 IN_M.n14 0.110917
R7902 IN_M.n50 IN_M.n49 0.110917
R7903 IN_M.n158 IN_M.n157 0.108833
R7904 IN_M.n48 IN_M.n47 0.108833
R7905 IN_M.n130 IN_M.n129 0.106502
R7906 IN_M.n20 IN_M.n19 0.106502
R7907 IN_M.n55 IN_M.n54 0.106502
R7908 IN_M.n195 IN_M.n194 0.106243
R7909 IN_M.n160 IN_M.n159 0.105998
R7910 IN_M.n85 IN_M.n84 0.105998
R7911 IN_M.n135 IN_M.n134 0.084875
R7912 IN_M.n142 IN_M.n141 0.084875
R7913 IN_M.n147 IN_M.n119 0.084875
R7914 IN_M.n163 IN_M.n162 0.084875
R7915 IN_M.n170 IN_M.n169 0.084875
R7916 IN_M.n177 IN_M.n176 0.084875
R7917 IN_M.n182 IN_M.n114 0.084875
R7918 IN_M.n189 IN_M.n113 0.084875
R7919 IN_M.n198 IN_M.n197 0.084875
R7920 IN_M.n205 IN_M.n204 0.084875
R7921 IN_M.n212 IN_M.n211 0.084875
R7922 IN_M.n102 IN_M.n101 0.084875
R7923 IN_M.n95 IN_M.n94 0.084875
R7924 IN_M.n88 IN_M.n87 0.084875
R7925 IN_M.n79 IN_M.n3 0.084875
R7926 IN_M.n72 IN_M.n4 0.084875
R7927 IN_M.n67 IN_M.n66 0.084875
R7928 IN_M.n60 IN_M.n59 0.084875
R7929 IN_M.n37 IN_M.n9 0.084875
R7930 IN_M.n32 IN_M.n31 0.084875
R7931 IN_M.n25 IN_M.n24 0.084875
R7932 IN_M.n126 IN_M.n122 0.0833125
R7933 IN_M.n51 IN_M.n7 0.0833125
R7934 IN_M.n16 IN_M.n12 0.0833125
R7935 IN_M.n140 IN_M.n120 0.08175
R7936 IN_M.n149 IN_M.n148 0.08175
R7937 IN_M.n156 IN_M.n155 0.08175
R7938 IN_M.n175 IN_M.n115 0.08175
R7939 IN_M.n184 IN_M.n183 0.08175
R7940 IN_M.n210 IN_M.n110 0.08175
R7941 IN_M.n100 IN_M.n0 0.08175
R7942 IN_M.n74 IN_M.n73 0.08175
R7943 IN_M.n65 IN_M.n5 0.08175
R7944 IN_M.n46 IN_M.n45 0.08175
R7945 IN_M.n39 IN_M.n38 0.08175
R7946 IN_M.n30 IN_M.n10 0.08175
R7947 IN_M.n154 IN_M.n118 0.078625
R7948 IN_M.n44 IN_M.n8 0.078625
R7949 IN_M.n133 IN_M.n121 0.0755
R7950 IN_M.n168 IN_M.n116 0.0755
R7951 IN_M.n191 IN_M.n190 0.0755
R7952 IN_M.n203 IN_M.n111 0.0755
R7953 IN_M.n93 IN_M.n1 0.0755
R7954 IN_M.n81 IN_M.n80 0.0755
R7955 IN_M.n58 IN_M.n6 0.0755
R7956 IN_M.n23 IN_M.n11 0.0755
R7957 IN_M.n128 IN_M.n127 0.06925
R7958 IN_M.n161 IN_M.n117 0.06925
R7959 IN_M.n196 IN_M.n112 0.06925
R7960 IN_M.n86 IN_M.n2 0.06925
R7961 IN_M.n53 IN_M.n52 0.06925
R7962 IN_M.n18 IN_M.n17 0.06925
R7963 IN_M.n106 IN_M.n105 0.0421667
R7964 IN_M.n216 IN_M.n215 0.0218477
R7965 IN_M.n128 IN_M.n126 0.016125
R7966 IN_M.n163 IN_M.n161 0.016125
R7967 IN_M.n198 IN_M.n196 0.016125
R7968 IN_M.n88 IN_M.n86 0.016125
R7969 IN_M.n53 IN_M.n51 0.016125
R7970 IN_M.n18 IN_M.n16 0.016125
R7971 IN_M.n219 IN_M.n216 0.0135011
R7972 IN_M.n109 IN_M.n106 0.0135011
R7973 IN_M.n135 IN_M.n133 0.009875
R7974 IN_M.n170 IN_M.n168 0.009875
R7975 IN_M.n191 IN_M.n189 0.009875
R7976 IN_M.n205 IN_M.n203 0.009875
R7977 IN_M.n95 IN_M.n93 0.009875
R7978 IN_M.n81 IN_M.n79 0.009875
R7979 IN_M.n60 IN_M.n58 0.009875
R7980 IN_M.n25 IN_M.n23 0.009875
R7981 IN_M.n156 IN_M.n154 0.00675
R7982 IN_M.n46 IN_M.n44 0.00675
R7983 IN_M.n218 IN_M.n217 0.00466667
R7984 IN_M.n108 IN_M.n107 0.00378079
R7985 IN_M.n142 IN_M.n140 0.003625
R7986 IN_M.n149 IN_M.n147 0.003625
R7987 IN_M.n177 IN_M.n175 0.003625
R7988 IN_M.n184 IN_M.n182 0.003625
R7989 IN_M.n212 IN_M.n210 0.003625
R7990 IN_M.n102 IN_M.n100 0.003625
R7991 IN_M.n74 IN_M.n72 0.003625
R7992 IN_M.n67 IN_M.n65 0.003625
R7993 IN_M.n39 IN_M.n37 0.003625
R7994 IN_M.n32 IN_M.n30 0.003625
R7995 IN_M.n219 IN_M.n218 0.00111601
R7996 IN_M.n109 IN_M.n108 0.00111601
R7997 IN_M.n213 IN_M.n212 0.000542675
R7998 IN_M.n206 IN_M.n205 0.000542675
R7999 IN_M.n199 IN_M.n198 0.000542675
R8000 IN_M.n189 IN_M.n188 0.000542675
R8001 IN_M.n182 IN_M.n181 0.000542675
R8002 IN_M.n178 IN_M.n177 0.000542675
R8003 IN_M.n171 IN_M.n170 0.000542675
R8004 IN_M.n164 IN_M.n163 0.000542675
R8005 IN_M.n157 IN_M.n156 0.000542675
R8006 IN_M.n147 IN_M.n146 0.000542675
R8007 IN_M.n143 IN_M.n142 0.000542675
R8008 IN_M.n136 IN_M.n135 0.000542675
R8009 IN_M.n126 IN_M.n125 0.000542675
R8010 IN_M.n16 IN_M.n15 0.000542675
R8011 IN_M.n26 IN_M.n25 0.000542675
R8012 IN_M.n33 IN_M.n32 0.000542675
R8013 IN_M.n37 IN_M.n36 0.000542675
R8014 IN_M.n47 IN_M.n46 0.000542675
R8015 IN_M.n51 IN_M.n50 0.000542675
R8016 IN_M.n61 IN_M.n60 0.000542675
R8017 IN_M.n68 IN_M.n67 0.000542675
R8018 IN_M.n72 IN_M.n71 0.000542675
R8019 IN_M.n79 IN_M.n78 0.000542675
R8020 IN_M.n89 IN_M.n88 0.000542675
R8021 IN_M.n96 IN_M.n95 0.000542675
R8022 IN_M.n103 IN_M.n102 0.000542675
R8023 IN_M.n154 IN_M.n153 0.000510684
R8024 IN_M.n44 IN_M.n43 0.000510684
R8025 IN_M.n129 IN_M.n128 0.000508707
R8026 IN_M.n133 IN_M.n132 0.000508707
R8027 IN_M.n140 IN_M.n139 0.000508707
R8028 IN_M.n150 IN_M.n149 0.000508707
R8029 IN_M.n161 IN_M.n160 0.000508707
R8030 IN_M.n168 IN_M.n167 0.000508707
R8031 IN_M.n175 IN_M.n174 0.000508707
R8032 IN_M.n185 IN_M.n184 0.000508707
R8033 IN_M.n192 IN_M.n191 0.000508707
R8034 IN_M.n196 IN_M.n195 0.000508707
R8035 IN_M.n203 IN_M.n202 0.000508707
R8036 IN_M.n210 IN_M.n209 0.000508707
R8037 IN_M.n100 IN_M.n99 0.000508707
R8038 IN_M.n93 IN_M.n92 0.000508707
R8039 IN_M.n86 IN_M.n85 0.000508707
R8040 IN_M.n82 IN_M.n81 0.000508707
R8041 IN_M.n75 IN_M.n74 0.000508707
R8042 IN_M.n65 IN_M.n64 0.000508707
R8043 IN_M.n58 IN_M.n57 0.000508707
R8044 IN_M.n54 IN_M.n53 0.000508707
R8045 IN_M.n40 IN_M.n39 0.000508707
R8046 IN_M.n30 IN_M.n29 0.000508707
R8047 IN_M.n23 IN_M.n22 0.000508707
R8048 IN_M.n19 IN_M.n18 0.000508707
R8049 a_46836_49340.n28 a_46836_49340.t47 8.53502
R8050 a_46836_49340.n30 a_46836_49340.t49 8.28993
R8051 a_46836_49340.n14 a_46836_49340.t30 7.5398
R8052 a_46836_49340.n0 a_46836_49340.t12 7.5398
R8053 a_46836_49340.t45 a_46836_49340.n49 6.90131
R8054 a_46836_49340.n49 a_46836_49340.t3 6.90131
R8055 a_46836_49340.n25 a_46836_49340.t37 6.90131
R8056 a_46836_49340.n11 a_46836_49340.t5 6.90131
R8057 a_46836_49340.n16 a_46836_49340.t32 6.83609
R8058 a_46836_49340.n2 a_46836_49340.t8 6.83609
R8059 a_46836_49340.n40 a_46836_49340.t6 6.83609
R8060 a_46836_49340.n40 a_46836_49340.t43 6.83609
R8061 a_46836_49340.n27 a_46836_49340.t34 6.82522
R8062 a_46836_49340.n13 a_46836_49340.t53 6.82522
R8063 a_46836_49340.n35 a_46836_49340.t56 6.82522
R8064 a_46836_49340.n35 a_46836_49340.t44 6.82522
R8065 a_46836_49340.n37 a_46836_49340.t1 6.81435
R8066 a_46836_49340.n37 a_46836_49340.t41 6.81435
R8067 a_46836_49340.n24 a_46836_49340.t28 6.80348
R8068 a_46836_49340.n10 a_46836_49340.t55 6.80348
R8069 a_46836_49340.n48 a_46836_49340.t61 6.80348
R8070 a_46836_49340.n48 a_46836_49340.t36 6.80348
R8071 a_46836_49340.n21 a_46836_49340.t38 6.78174
R8072 a_46836_49340.n7 a_46836_49340.t4 6.78174
R8073 a_46836_49340.n45 a_46836_49340.t2 6.78174
R8074 a_46836_49340.n45 a_46836_49340.t16 6.78174
R8075 a_46836_49340.n18 a_46836_49340.t23 6.76001
R8076 a_46836_49340.n4 a_46836_49340.t63 6.76001
R8077 a_46836_49340.n42 a_46836_49340.t52 6.76001
R8078 a_46836_49340.n42 a_46836_49340.t29 6.76001
R8079 a_46836_49340.n15 a_46836_49340.t31 6.73827
R8080 a_46836_49340.n1 a_46836_49340.t9 6.73827
R8081 a_46836_49340.n39 a_46836_49340.t7 6.73827
R8082 a_46836_49340.n39 a_46836_49340.t42 6.73827
R8083 a_46836_49340.n26 a_46836_49340.t26 6.7274
R8084 a_46836_49340.n12 a_46836_49340.t62 6.7274
R8085 a_46836_49340.n36 a_46836_49340.t15 6.7274
R8086 a_46836_49340.n36 a_46836_49340.t33 6.7274
R8087 a_46836_49340.n23 a_46836_49340.t27 6.70566
R8088 a_46836_49340.n9 a_46836_49340.t10 6.70566
R8089 a_46836_49340.n47 a_46836_49340.t14 6.70566
R8090 a_46836_49340.n47 a_46836_49340.t35 6.70566
R8091 a_46836_49340.n20 a_46836_49340.t20 6.68392
R8092 a_46836_49340.n6 a_46836_49340.t0 6.68392
R8093 a_46836_49340.n44 a_46836_49340.t54 6.68392
R8094 a_46836_49340.n44 a_46836_49340.t24 6.68392
R8095 a_46836_49340.n17 a_46836_49340.t39 6.66218
R8096 a_46836_49340.n3 a_46836_49340.t65 6.66218
R8097 a_46836_49340.n14 a_46836_49340.t21 6.64044
R8098 a_46836_49340.n0 a_46836_49340.t57 6.64044
R8099 a_46836_49340.n38 a_46836_49340.t13 6.64044
R8100 a_46836_49340.n38 a_46836_49340.t25 6.64044
R8101 a_46836_49340.n22 a_46836_49340.t17 6.60783
R8102 a_46836_49340.n8 a_46836_49340.t60 6.60783
R8103 a_46836_49340.n41 a_46836_49340.t59 6.60783
R8104 a_46836_49340.n41 a_46836_49340.t18 6.60783
R8105 a_46836_49340.n46 a_46836_49340.t11 6.60783
R8106 a_46836_49340.n46 a_46836_49340.t22 6.60783
R8107 a_46836_49340.n19 a_46836_49340.t40 6.58609
R8108 a_46836_49340.n5 a_46836_49340.t64 6.58609
R8109 a_46836_49340.n43 a_46836_49340.t58 6.58609
R8110 a_46836_49340.n43 a_46836_49340.t19 6.58609
R8111 a_46836_49340.n33 a_46836_49340.n32 5.88188
R8112 a_46836_49340.n29 a_46836_49340.t50 5.72994
R8113 a_46836_49340.n31 a_46836_49340.t46 5.72994
R8114 a_46836_49340.n28 a_46836_49340.t48 5.71419
R8115 a_46836_49340.n30 a_46836_49340.t51 5.71419
R8116 a_46836_49340.n29 a_46836_49340.n28 2.38339
R8117 a_46836_49340.n31 a_46836_49340.n30 2.32334
R8118 a_46836_49340.n34 a_46836_49340.n13 2.21875
R8119 a_46836_49340.n33 a_46836_49340.n27 1.93029
R8120 a_46836_49340.n35 a_46836_49340.n34 1.93029
R8121 a_46836_49340.n32 a_46836_49340.n29 1.07166
R8122 a_46836_49340.n41 a_46836_49340.n40 0.737107
R8123 a_46836_49340.n26 a_46836_49340.n25 0.725946
R8124 a_46836_49340.n22 a_46836_49340.n21 0.725946
R8125 a_46836_49340.n19 a_46836_49340.n18 0.725946
R8126 a_46836_49340.n17 a_46836_49340.n16 0.725946
R8127 a_46836_49340.n12 a_46836_49340.n11 0.725946
R8128 a_46836_49340.n8 a_46836_49340.n7 0.725946
R8129 a_46836_49340.n5 a_46836_49340.n4 0.725946
R8130 a_46836_49340.n3 a_46836_49340.n2 0.725946
R8131 a_46836_49340.n49 a_46836_49340.n36 0.725946
R8132 a_46836_49340.n46 a_46836_49340.n45 0.725946
R8133 a_46836_49340.n43 a_46836_49340.n42 0.725946
R8134 a_46836_49340.n38 a_46836_49340.n37 0.725946
R8135 a_46836_49340.n27 a_46836_49340.n26 0.670143
R8136 a_46836_49340.n25 a_46836_49340.n24 0.670143
R8137 a_46836_49340.n24 a_46836_49340.n23 0.670143
R8138 a_46836_49340.n23 a_46836_49340.n22 0.670143
R8139 a_46836_49340.n21 a_46836_49340.n20 0.670143
R8140 a_46836_49340.n20 a_46836_49340.n19 0.670143
R8141 a_46836_49340.n18 a_46836_49340.n17 0.670143
R8142 a_46836_49340.n16 a_46836_49340.n15 0.670143
R8143 a_46836_49340.n15 a_46836_49340.n14 0.670143
R8144 a_46836_49340.n13 a_46836_49340.n12 0.670143
R8145 a_46836_49340.n11 a_46836_49340.n10 0.670143
R8146 a_46836_49340.n10 a_46836_49340.n9 0.670143
R8147 a_46836_49340.n9 a_46836_49340.n8 0.670143
R8148 a_46836_49340.n7 a_46836_49340.n6 0.670143
R8149 a_46836_49340.n6 a_46836_49340.n5 0.670143
R8150 a_46836_49340.n4 a_46836_49340.n3 0.670143
R8151 a_46836_49340.n2 a_46836_49340.n1 0.670143
R8152 a_46836_49340.n1 a_46836_49340.n0 0.670143
R8153 a_46836_49340.n36 a_46836_49340.n35 0.670143
R8154 a_46836_49340.n49 a_46836_49340.n48 0.670143
R8155 a_46836_49340.n48 a_46836_49340.n47 0.670143
R8156 a_46836_49340.n47 a_46836_49340.n46 0.670143
R8157 a_46836_49340.n45 a_46836_49340.n44 0.670143
R8158 a_46836_49340.n44 a_46836_49340.n43 0.670143
R8159 a_46836_49340.n40 a_46836_49340.n39 0.670143
R8160 a_46836_49340.n39 a_46836_49340.n38 0.670143
R8161 a_46836_49340.n42 a_46836_49340.n41 0.658982
R8162 a_46836_49340.n34 a_46836_49340.n33 0.288962
R8163 a_46836_49340.n32 a_46836_49340.n31 0.121657
R8164 IN_P.n217 IN_P.t15 746.848
R8165 IN_P.n11 IN_P.t23 746.846
R8166 IN_P.n10 IN_P.t1 746.846
R8167 IN_P.n9 IN_P.t2 746.846
R8168 IN_P.n8 IN_P.t16 746.846
R8169 IN_P.n7 IN_P.t22 746.846
R8170 IN_P.n6 IN_P.t14 746.846
R8171 IN_P.n5 IN_P.t20 746.846
R8172 IN_P.n4 IN_P.t5 746.846
R8173 IN_P.n3 IN_P.t21 746.846
R8174 IN_P.n2 IN_P.t26 746.846
R8175 IN_P.n1 IN_P.t27 746.846
R8176 IN_P.n0 IN_P.t11 746.846
R8177 IN_P.n107 IN_P.t28 746.846
R8178 IN_P.n110 IN_P.t29 746.846
R8179 IN_P.n111 IN_P.t13 746.846
R8180 IN_P.n112 IN_P.t12 746.846
R8181 IN_P.n113 IN_P.t7 746.846
R8182 IN_P.n114 IN_P.t24 746.846
R8183 IN_P.n115 IN_P.t6 746.846
R8184 IN_P.n116 IN_P.t0 746.846
R8185 IN_P.n117 IN_P.t8 746.846
R8186 IN_P.n118 IN_P.t3 746.846
R8187 IN_P.n119 IN_P.t18 746.846
R8188 IN_P.n120 IN_P.t17 746.846
R8189 IN_P.n121 IN_P.t9 746.846
R8190 IN_P.n122 IN_P.t19 746.309
R8191 IN_P.n12 IN_P.t4 746.309
R8192 IN_P.n123 IN_P.t10 374.077
R8193 IN_P.n13 IN_P.t25 374.077
R8194 IN_P IN_P.n220 4.62423
R8195 IN_P.n220 IN_P.n109 2.85474
R8196 IN_P.n220 IN_P.n219 2.83326
R8197 IN_P.n124 IN_P.n123 2.43766
R8198 IN_P.n14 IN_P.n13 2.43766
R8199 IN_P.n159 IN_P.n158 2.34135
R8200 IN_P.n49 IN_P.n48 2.34135
R8201 IN_P.n166 IN_P.n165 2.33827
R8202 IN_P.n201 IN_P.n200 2.33827
R8203 IN_P.n56 IN_P.n55 2.33827
R8204 IN_P.n91 IN_P.n90 2.33827
R8205 IN_P.n42 IN_P.n41 2.33055
R8206 IN_P.n145 IN_P.n144 2.32981
R8207 IN_P.n180 IN_P.n179 2.32981
R8208 IN_P.n35 IN_P.n34 2.32981
R8209 IN_P.n70 IN_P.n69 2.32981
R8210 IN_P.n138 IN_P.n137 2.32981
R8211 IN_P.n173 IN_P.n172 2.32981
R8212 IN_P.n208 IN_P.n207 2.32981
R8213 IN_P.n28 IN_P.n27 2.32981
R8214 IN_P.n63 IN_P.n62 2.32981
R8215 IN_P.n98 IN_P.n97 2.32981
R8216 IN_P.n152 IN_P.n151 2.3298
R8217 IN_P.n187 IN_P.n186 2.3298
R8218 IN_P.n77 IN_P.n76 2.3298
R8219 IN_P.n84 IN_P.n83 2.32516
R8220 IN_P.n194 IN_P.n193 2.32442
R8221 IN_P.n131 IN_P.n130 2.32441
R8222 IN_P.n21 IN_P.n20 2.32441
R8223 IN_P.n105 IN_P.n104 2.31935
R8224 IN_P.n215 IN_P.n214 2.29822
R8225 IN_P.n144 IN_P.n143 0.1243
R8226 IN_P.n179 IN_P.n178 0.1243
R8227 IN_P.n214 IN_P.n213 0.1243
R8228 IN_P.n34 IN_P.n33 0.1243
R8229 IN_P.n69 IN_P.n68 0.1243
R8230 IN_P.n104 IN_P.n103 0.1243
R8231 IN_P.n146 IN_P.n145 0.123792
R8232 IN_P.n181 IN_P.n180 0.123792
R8233 IN_P.n36 IN_P.n35 0.123792
R8234 IN_P.n71 IN_P.n70 0.123792
R8235 IN_P.n137 IN_P.n136 0.123283
R8236 IN_P.n172 IN_P.n171 0.123283
R8237 IN_P.n207 IN_P.n206 0.123283
R8238 IN_P.n27 IN_P.n26 0.123283
R8239 IN_P.n62 IN_P.n61 0.123283
R8240 IN_P.n97 IN_P.n96 0.123283
R8241 IN_P.n188 IN_P.n187 0.122774
R8242 IN_P.n78 IN_P.n77 0.122774
R8243 IN_P.n151 IN_P.n150 0.121147
R8244 IN_P.n186 IN_P.n185 0.121147
R8245 IN_P.n41 IN_P.n40 0.121147
R8246 IN_P.n76 IN_P.n75 0.121147
R8247 IN_P.n139 IN_P.n138 0.120641
R8248 IN_P.n174 IN_P.n173 0.120641
R8249 IN_P.n209 IN_P.n208 0.120641
R8250 IN_P.n29 IN_P.n28 0.120641
R8251 IN_P.n64 IN_P.n63 0.120641
R8252 IN_P.n99 IN_P.n98 0.120641
R8253 IN_P.n43 IN_P.n42 0.114687
R8254 IN_P.n153 IN_P.n152 0.11444
R8255 IN_P.n193 IN_P.n192 0.113826
R8256 IN_P.n83 IN_P.n82 0.113826
R8257 IN_P.n132 IN_P.n131 0.11332
R8258 IN_P.n167 IN_P.n166 0.11332
R8259 IN_P.n202 IN_P.n201 0.11332
R8260 IN_P.n22 IN_P.n21 0.11332
R8261 IN_P.n57 IN_P.n56 0.11332
R8262 IN_P.n92 IN_P.n91 0.11332
R8263 IN_P.n165 IN_P.n164 0.113
R8264 IN_P.n200 IN_P.n199 0.113
R8265 IN_P.n55 IN_P.n54 0.113
R8266 IN_P.n90 IN_P.n89 0.113
R8267 IN_P.n125 IN_P.n124 0.110917
R8268 IN_P.n15 IN_P.n14 0.110917
R8269 IN_P.n158 IN_P.n157 0.108833
R8270 IN_P.n48 IN_P.n47 0.108833
R8271 IN_P.n130 IN_P.n129 0.106502
R8272 IN_P.n20 IN_P.n19 0.106502
R8273 IN_P.n85 IN_P.n84 0.106243
R8274 IN_P.n160 IN_P.n159 0.105998
R8275 IN_P.n195 IN_P.n194 0.105998
R8276 IN_P.n50 IN_P.n49 0.105998
R8277 IN_P.n212 IN_P.n211 0.084875
R8278 IN_P.n205 IN_P.n204 0.084875
R8279 IN_P.n198 IN_P.n197 0.084875
R8280 IN_P.n189 IN_P.n113 0.084875
R8281 IN_P.n182 IN_P.n114 0.084875
R8282 IN_P.n177 IN_P.n176 0.084875
R8283 IN_P.n170 IN_P.n169 0.084875
R8284 IN_P.n163 IN_P.n162 0.084875
R8285 IN_P.n147 IN_P.n119 0.084875
R8286 IN_P.n142 IN_P.n141 0.084875
R8287 IN_P.n135 IN_P.n134 0.084875
R8288 IN_P.n25 IN_P.n24 0.084875
R8289 IN_P.n32 IN_P.n31 0.084875
R8290 IN_P.n37 IN_P.n9 0.084875
R8291 IN_P.n53 IN_P.n52 0.084875
R8292 IN_P.n60 IN_P.n59 0.084875
R8293 IN_P.n67 IN_P.n66 0.084875
R8294 IN_P.n72 IN_P.n4 0.084875
R8295 IN_P.n79 IN_P.n3 0.084875
R8296 IN_P.n88 IN_P.n87 0.084875
R8297 IN_P.n95 IN_P.n94 0.084875
R8298 IN_P.n102 IN_P.n101 0.084875
R8299 IN_P.n126 IN_P.n122 0.0833125
R8300 IN_P.n16 IN_P.n12 0.0833125
R8301 IN_P.n210 IN_P.n110 0.08175
R8302 IN_P.n184 IN_P.n183 0.08175
R8303 IN_P.n175 IN_P.n115 0.08175
R8304 IN_P.n156 IN_P.n155 0.08175
R8305 IN_P.n149 IN_P.n148 0.08175
R8306 IN_P.n140 IN_P.n120 0.08175
R8307 IN_P.n30 IN_P.n10 0.08175
R8308 IN_P.n39 IN_P.n38 0.08175
R8309 IN_P.n46 IN_P.n45 0.08175
R8310 IN_P.n65 IN_P.n5 0.08175
R8311 IN_P.n74 IN_P.n73 0.08175
R8312 IN_P.n100 IN_P.n0 0.08175
R8313 IN_P.n154 IN_P.n118 0.078625
R8314 IN_P.n44 IN_P.n8 0.078625
R8315 IN_P.n203 IN_P.n111 0.0755
R8316 IN_P.n191 IN_P.n190 0.0755
R8317 IN_P.n168 IN_P.n116 0.0755
R8318 IN_P.n133 IN_P.n121 0.0755
R8319 IN_P.n23 IN_P.n11 0.0755
R8320 IN_P.n58 IN_P.n6 0.0755
R8321 IN_P.n81 IN_P.n80 0.0755
R8322 IN_P.n93 IN_P.n1 0.0755
R8323 IN_P.n196 IN_P.n112 0.06925
R8324 IN_P.n161 IN_P.n117 0.06925
R8325 IN_P.n128 IN_P.n127 0.06925
R8326 IN_P.n18 IN_P.n17 0.06925
R8327 IN_P.n51 IN_P.n7 0.06925
R8328 IN_P.n86 IN_P.n2 0.06925
R8329 IN_P.n216 IN_P.n215 0.0421667
R8330 IN_P.n106 IN_P.n105 0.0218477
R8331 IN_P.n198 IN_P.n196 0.016125
R8332 IN_P.n163 IN_P.n161 0.016125
R8333 IN_P.n128 IN_P.n126 0.016125
R8334 IN_P.n18 IN_P.n16 0.016125
R8335 IN_P.n53 IN_P.n51 0.016125
R8336 IN_P.n88 IN_P.n86 0.016125
R8337 IN_P.n219 IN_P.n216 0.0135011
R8338 IN_P.n109 IN_P.n106 0.0135011
R8339 IN_P.n205 IN_P.n203 0.009875
R8340 IN_P.n191 IN_P.n189 0.009875
R8341 IN_P.n170 IN_P.n168 0.009875
R8342 IN_P.n135 IN_P.n133 0.009875
R8343 IN_P.n25 IN_P.n23 0.009875
R8344 IN_P.n60 IN_P.n58 0.009875
R8345 IN_P.n81 IN_P.n79 0.009875
R8346 IN_P.n95 IN_P.n93 0.009875
R8347 IN_P.n156 IN_P.n154 0.00675
R8348 IN_P.n46 IN_P.n44 0.00675
R8349 IN_P.n108 IN_P.n107 0.00466667
R8350 IN_P.n218 IN_P.n217 0.00378079
R8351 IN_P.n212 IN_P.n210 0.003625
R8352 IN_P.n184 IN_P.n182 0.003625
R8353 IN_P.n177 IN_P.n175 0.003625
R8354 IN_P.n149 IN_P.n147 0.003625
R8355 IN_P.n142 IN_P.n140 0.003625
R8356 IN_P.n32 IN_P.n30 0.003625
R8357 IN_P.n39 IN_P.n37 0.003625
R8358 IN_P.n67 IN_P.n65 0.003625
R8359 IN_P.n74 IN_P.n72 0.003625
R8360 IN_P.n102 IN_P.n100 0.003625
R8361 IN_P.n219 IN_P.n218 0.00111601
R8362 IN_P.n109 IN_P.n108 0.00111601
R8363 IN_P.n126 IN_P.n125 0.000542675
R8364 IN_P.n136 IN_P.n135 0.000542675
R8365 IN_P.n143 IN_P.n142 0.000542675
R8366 IN_P.n147 IN_P.n146 0.000542675
R8367 IN_P.n157 IN_P.n156 0.000542675
R8368 IN_P.n164 IN_P.n163 0.000542675
R8369 IN_P.n171 IN_P.n170 0.000542675
R8370 IN_P.n178 IN_P.n177 0.000542675
R8371 IN_P.n182 IN_P.n181 0.000542675
R8372 IN_P.n189 IN_P.n188 0.000542675
R8373 IN_P.n199 IN_P.n198 0.000542675
R8374 IN_P.n206 IN_P.n205 0.000542675
R8375 IN_P.n213 IN_P.n212 0.000542675
R8376 IN_P.n103 IN_P.n102 0.000542675
R8377 IN_P.n96 IN_P.n95 0.000542675
R8378 IN_P.n89 IN_P.n88 0.000542675
R8379 IN_P.n79 IN_P.n78 0.000542675
R8380 IN_P.n72 IN_P.n71 0.000542675
R8381 IN_P.n68 IN_P.n67 0.000542675
R8382 IN_P.n61 IN_P.n60 0.000542675
R8383 IN_P.n54 IN_P.n53 0.000542675
R8384 IN_P.n47 IN_P.n46 0.000542675
R8385 IN_P.n37 IN_P.n36 0.000542675
R8386 IN_P.n33 IN_P.n32 0.000542675
R8387 IN_P.n26 IN_P.n25 0.000542675
R8388 IN_P.n16 IN_P.n15 0.000542675
R8389 IN_P.n154 IN_P.n153 0.000510684
R8390 IN_P.n44 IN_P.n43 0.000510684
R8391 IN_P.n210 IN_P.n209 0.000508707
R8392 IN_P.n203 IN_P.n202 0.000508707
R8393 IN_P.n196 IN_P.n195 0.000508707
R8394 IN_P.n192 IN_P.n191 0.000508707
R8395 IN_P.n185 IN_P.n184 0.000508707
R8396 IN_P.n175 IN_P.n174 0.000508707
R8397 IN_P.n168 IN_P.n167 0.000508707
R8398 IN_P.n161 IN_P.n160 0.000508707
R8399 IN_P.n150 IN_P.n149 0.000508707
R8400 IN_P.n140 IN_P.n139 0.000508707
R8401 IN_P.n133 IN_P.n132 0.000508707
R8402 IN_P.n129 IN_P.n128 0.000508707
R8403 IN_P.n19 IN_P.n18 0.000508707
R8404 IN_P.n23 IN_P.n22 0.000508707
R8405 IN_P.n30 IN_P.n29 0.000508707
R8406 IN_P.n40 IN_P.n39 0.000508707
R8407 IN_P.n51 IN_P.n50 0.000508707
R8408 IN_P.n58 IN_P.n57 0.000508707
R8409 IN_P.n65 IN_P.n64 0.000508707
R8410 IN_P.n75 IN_P.n74 0.000508707
R8411 IN_P.n82 IN_P.n81 0.000508707
R8412 IN_P.n86 IN_P.n85 0.000508707
R8413 IN_P.n93 IN_P.n92 0.000508707
R8414 IN_P.n100 IN_P.n99 0.000508707
R8415 bias21.n22 bias21.t38 65.7944
R8416 bias21 bias21.n14 40.7763
R8417 bias21.n15 bias21.t4 22.674
R8418 bias21.n17 bias21.t6 21.4485
R8419 bias21.n16 bias21.t0 21.4435
R8420 bias21.n15 bias21.t2 21.4435
R8421 bias21.n18 bias21.t5 15.0848
R8422 bias21.n20 bias21.t7 13.9238
R8423 bias21.n19 bias21.t1 13.9238
R8424 bias21.n18 bias21.t3 13.9238
R8425 bias21.n12 bias21.t14 6.90131
R8426 bias21.n12 bias21.t28 6.90131
R8427 bias21.n3 bias21.t11 6.83609
R8428 bias21.n3 bias21.t25 6.83609
R8429 bias21.n14 bias21.t12 6.82522
R8430 bias21.n14 bias21.t27 6.82522
R8431 bias21.n0 bias21.t9 6.81435
R8432 bias21.n0 bias21.t22 6.81435
R8433 bias21.n11 bias21.t36 6.80348
R8434 bias21.n11 bias21.t20 6.80348
R8435 bias21.n8 bias21.t15 6.78174
R8436 bias21.n8 bias21.t29 6.78174
R8437 bias21.n5 bias21.t32 6.76001
R8438 bias21.n5 bias21.t13 6.76001
R8439 bias21.n2 bias21.t10 6.73827
R8440 bias21.n2 bias21.t24 6.73827
R8441 bias21.n13 bias21.t33 6.7274
R8442 bias21.n13 bias21.t18 6.7274
R8443 bias21.n10 bias21.t35 6.70566
R8444 bias21.n10 bias21.t19 6.70566
R8445 bias21.n7 bias21.t23 6.68392
R8446 bias21.n7 bias21.t37 6.68392
R8447 bias21.n1 bias21.t26 6.64044
R8448 bias21.n1 bias21.t8 6.64044
R8449 bias21.n4 bias21.t16 6.60783
R8450 bias21.n4 bias21.t30 6.60783
R8451 bias21.n9 bias21.t21 6.60783
R8452 bias21.n9 bias21.t34 6.60783
R8453 bias21.n6 bias21.t17 6.58609
R8454 bias21.n6 bias21.t31 6.58609
R8455 bias21 bias21.n22 3.18783
R8456 bias21.n22 bias21.n21 2.90116
R8457 bias21.n16 bias21.n15 1.231
R8458 bias21.n17 bias21.n16 1.22365
R8459 bias21.n19 bias21.n18 1.16148
R8460 bias21.n20 bias21.n19 1.16148
R8461 bias21.n21 bias21.n17 0.898924
R8462 bias21.n4 bias21.n3 0.737107
R8463 bias21.n13 bias21.n12 0.725946
R8464 bias21.n9 bias21.n8 0.725946
R8465 bias21.n6 bias21.n5 0.725946
R8466 bias21.n1 bias21.n0 0.725946
R8467 bias21.n14 bias21.n13 0.670143
R8468 bias21.n12 bias21.n11 0.670143
R8469 bias21.n11 bias21.n10 0.670143
R8470 bias21.n10 bias21.n9 0.670143
R8471 bias21.n8 bias21.n7 0.670143
R8472 bias21.n7 bias21.n6 0.670143
R8473 bias21.n3 bias21.n2 0.670143
R8474 bias21.n2 bias21.n1 0.670143
R8475 bias21.n5 bias21.n4 0.658982
R8476 bias21.n21 bias21.n20 0.402867
R8477 m11m12 m11m12.t30 13.1423
R8478 m11m12.n28 m11m12.n13 12.4583
R8479 m11m12.n28 m11m12.n27 6.07595
R8480 m11m12.n0 m11m12.t28 4.44742
R8481 m11m12.n14 m11m12.t6 4.42883
R8482 m11m12 m11m12.n28 3.55758
R8483 m11m12.n17 m11m12.t29 3.48118
R8484 m11m12.n18 m11m12.t4 3.48118
R8485 m11m12.n19 m11m12.t17 3.48118
R8486 m11m12.n20 m11m12.t15 3.48118
R8487 m11m12.n21 m11m12.t13 3.48118
R8488 m11m12.n22 m11m12.t10 3.48118
R8489 m11m12.n23 m11m12.t19 3.48118
R8490 m11m12.n24 m11m12.t24 3.48118
R8491 m11m12.n25 m11m12.t22 3.48118
R8492 m11m12.n26 m11m12.t20 3.48118
R8493 m11m12.n27 m11m12.t2 3.48118
R8494 m11m12.n13 m11m12.t25 3.48118
R8495 m11m12.n12 m11m12.t12 3.48118
R8496 m11m12.n11 m11m12.t14 3.48118
R8497 m11m12.n10 m11m12.t16 3.48118
R8498 m11m12.n9 m11m12.t11 3.48118
R8499 m11m12.n8 m11m12.t5 3.48118
R8500 m11m12.n7 m11m12.t7 3.48118
R8501 m11m12.n6 m11m12.t8 3.48118
R8502 m11m12.n5 m11m12.t9 3.48118
R8503 m11m12.n4 m11m12.t27 3.48118
R8504 m11m12.n3 m11m12.t18 3.48118
R8505 m11m12.n2 m11m12.t21 3.48118
R8506 m11m12.n1 m11m12.t23 3.48118
R8507 m11m12.n0 m11m12.t26 3.48118
R8508 m11m12.n16 m11m12.t0 3.48118
R8509 m11m12.n15 m11m12.t1 3.48118
R8510 m11m12.n14 m11m12.t3 3.48118
R8511 m11m12.n1 m11m12.n0 0.966748
R8512 m11m12.n2 m11m12.n1 0.966748
R8513 m11m12.n3 m11m12.n2 0.966748
R8514 m11m12.n4 m11m12.n3 0.966748
R8515 m11m12.n5 m11m12.n4 0.966748
R8516 m11m12.n6 m11m12.n5 0.966748
R8517 m11m12.n7 m11m12.n6 0.966748
R8518 m11m12.n8 m11m12.n7 0.966748
R8519 m11m12.n9 m11m12.n8 0.966748
R8520 m11m12.n10 m11m12.n9 0.966748
R8521 m11m12.n11 m11m12.n10 0.966748
R8522 m11m12.n12 m11m12.n11 0.966748
R8523 m11m12.n13 m11m12.n12 0.966748
R8524 m11m12.n27 m11m12.n26 0.948155
R8525 m11m12.n26 m11m12.n25 0.948155
R8526 m11m12.n25 m11m12.n24 0.948155
R8527 m11m12.n24 m11m12.n23 0.948155
R8528 m11m12.n23 m11m12.n22 0.948155
R8529 m11m12.n22 m11m12.n21 0.948155
R8530 m11m12.n21 m11m12.n20 0.948155
R8531 m11m12.n20 m11m12.n19 0.948155
R8532 m11m12.n19 m11m12.n18 0.948155
R8533 m11m12.n18 m11m12.n17 0.948155
R8534 m11m12.n15 m11m12.n14 0.948155
R8535 m11m12.n16 m11m12.n15 0.948155
R8536 m11m12.n17 m11m12.n16 0.948155
C0 m1m2 VB_A 12.1f
C1 m1m2 dummy_9 30.6f
C2 dummy_4 bias21 0.406f
C3 bias3 m3m4 1.4f
C4 dummy_2 m9m10 2.69f
C5 bias1 m1m2 0.172p
C6 bias3 OUT 0.978f
C7 bias3 m11m12 0.374f
C8 dummy_4 m3m4 1.44f
C9 dummy_3 bias21 0.963f
C10 dummy_2 m1m2 2.65f
C11 IN_M IN_P 3.48f
C12 dummy_3 VB_B 50.4f
C13 bias3 VB_A 0.978f
C14 bias21 VCC 98.6f
C15 dummy_100 IB 24.6f
C16 dummy_3 m3m4 2.84f
C17 dummy_4 m11m12 1.08f
C18 m9m10 m1m2 99f
C19 VCC VB_B 0.923f
C20 bias3 IB 0.978f
C21 bias21 VB_B 1.01f
C22 dummy_3 OUT 2.64f
C23 bias3 m1_49040_35916# 0.406f
C24 bias21 m3m4 0.0154f
C25 dummy_3 m11m12 20.7f
C26 VCC OUT 11.1f
C27 bias21 OUT 0.978f
C28 bias3 IN_M 11.7f
C29 m3m4 VB_B 12.8f
C30 dummy_3 bias1 1.43f
C31 bias21 m11m12 0.948f
C32 VCC VB_A 94.8f
C33 VB_B OUT 11.7f
C34 dummy_9 VCC 0.285p
C35 m11m12 VB_B 12.6f
C36 m3m4 OUT 18.9f
C37 bias21 VB_A 1f
C38 bias1 VCC 3.16p
C39 m3m4 m11m12 0.403f
C40 VCC IB 40.3f
C41 m1_49040_35916# VCC 1.83f
C42 bias1 VB_B 11.2f
C43 dummy_2 VCC 17.3f
C44 m11m12 OUT 0.733f
C45 bias21 IB 1.01f
C46 bias21 m1_49040_35916# 0.27f
C47 bias21 dummy_2 0.89f
C48 m3m4 bias1 0.733f
C49 VCC IN_M 17.1f
C50 OUT VB_A 12.7f
C51 m9m10 VCC 0.435p
C52 bias1 OUT 1.61f
C53 VCC IN_P 15.8f
C54 bias21 IN_P 11.8f
C55 bias1 VB_A 13.2f
C56 m1m2 VCC 0.441p
C57 dummy_2 OUT 15.7f
C58 bias1 dummy_9 0.205p
C59 bias3 dummy_4 9.83f
C60 m9m10 OUT 0.738f
C61 dummy_2 VB_A 50.4f
C62 dummy_100 VCC 13.8f
C63 bias1 dummy_2 2.5f
C64 bias3 VCC 0.102p
C65 m9m10 VB_A 11.7f
C66 m9m10 dummy_9 31.1f
C67 bias3 bias21 10.1f
C68 bias1 m9m10 0.189p
C69 bias3 VB_B 0.978f
.ends

